-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

--library UNISIM;
--	use UNISIM.Vcomponents.all;

entity rom_oa is
port (
	CLK  : in  std_logic;
	ADDR : in  std_logic_vector(13 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of rom_oa is


	type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"4C",x"CC",x"EC",x"4C",x"71",x"C4",x"72",x"C9", -- 0x0000
		x"91",x"C6",x"86",x"E9",x"D0",x"E9",x"15",x"CD", -- 0x0008
		x"18",x"CD",x"11",x"CA",x"50",x"DA",x"A0",x"DA", -- 0x0010
		x"DD",x"D9",x"66",x"D9",x"84",x"DA",x"A0",x"DA", -- 0x0018
		x"54",x"C8",x"FC",x"C7",x"08",x"C8",x"97",x"CE", -- 0x0020
		x"3B",x"CA",x"54",x"CD",x"7D",x"D1",x"CD",x"CC", -- 0x0028
		x"88",x"CD",x"1B",x"CB",x"E4",x"C9",x"BC",x"C9", -- 0x0030
		x"6F",x"CA",x"51",x"C9",x"C7",x"C9",x"11",x"CA", -- 0x0038
		x"98",x"CA",x"CD",x"EB",x"E6",x"EB",x"0B",x"EC", -- 0x0040
		x"20",x"EC",x"32",x"EC",x"B4",x"FA",x"CA",x"FA", -- 0x0048
		x"E0",x"FA",x"9E",x"FA",x"FB",x"EA",x"FB",x"EA", -- 0x0050
		x"FB",x"EA",x"EF",x"EA",x"EF",x"EA",x"EF",x"EA", -- 0x0058
		x"EF",x"EA",x"EF",x"EA",x"EF",x"EA",x"EF",x"EA", -- 0x0060
		x"FB",x"EA",x"FB",x"EA",x"70",x"C9",x"C1",x"CA", -- 0x0068
		x"57",x"D9",x"5A",x"E8",x"08",x"E9",x"B9",x"D4", -- 0x0070
		x"4E",x"D9",x"AA",x"CB",x"9F",x"C9",x"47",x"C7", -- 0x0078
		x"0C",x"C7",x"45",x"CD",x"45",x"E9",x"12",x"CD", -- 0x0080
		x"ED",x"C6",x"21",x"DF",x"BD",x"DF",x"49",x"DF", -- 0x0088
		x"21",x"00",x"7E",x"D4",x"A6",x"D4",x"B5",x"D9", -- 0x0090
		x"FB",x"02",x"2E",x"E2",x"4F",x"E3",x"AF",x"DC", -- 0x0098
		x"AA",x"E2",x"8B",x"E3",x"92",x"E3",x"DB",x"E3", -- 0x00A0
		x"3F",x"E4",x"38",x"D9",x"83",x"D9",x"D4",x"DD", -- 0x00A8
		x"A6",x"D8",x"93",x"D5",x"D7",x"D8",x"B5",x"D8", -- 0x00B0
		x"16",x"D8",x"77",x"DE",x"0F",x"DF",x"0B",x"DF", -- 0x00B8
		x"DA",x"DA",x"3F",x"DA",x"45",x"EC",x"2A",x"D8", -- 0x00C0
		x"56",x"D8",x"61",x"D8",x"79",x"24",x"DB",x"79", -- 0x00C8
		x"0D",x"DB",x"7B",x"EF",x"DC",x"7B",x"E6",x"DD", -- 0x00D0
		x"7F",x"37",x"E2",x"50",x"E5",x"D0",x"46",x"E2", -- 0x00D8
		x"D0",x"7D",x"70",x"E2",x"5A",x"3B",x"D0",x"64", -- 0x00E0
		x"12",x"D1",x"45",x"4E",x"C4",x"45",x"44",x"49", -- 0x00E8
		x"D4",x"53",x"54",x"4F",x"52",x"C5",x"52",x"45", -- 0x00F0
		x"43",x"41",x"4C",x"CC",x"54",x"52",x"4F",x"CE", -- 0x00F8
		x"54",x"52",x"4F",x"46",x"C6",x"50",x"4F",x"D0", -- 0x0100
		x"50",x"4C",x"4F",x"D4",x"50",x"55",x"4C",x"CC", -- 0x0108
		x"4C",x"4F",x"52",x"45",x"D3",x"44",x"4F",x"4B", -- 0x0110
		x"C5",x"52",x"45",x"50",x"45",x"41",x"D4",x"55", -- 0x0118
		x"4E",x"54",x"49",x"CC",x"46",x"4F",x"D2",x"4C", -- 0x0120
		x"4C",x"49",x"53",x"D4",x"4C",x"50",x"52",x"49", -- 0x0128
		x"4E",x"D4",x"4E",x"45",x"58",x"D4",x"44",x"41", -- 0x0130
		x"54",x"C1",x"49",x"4E",x"50",x"55",x"D4",x"44", -- 0x0138
		x"49",x"CD",x"43",x"4C",x"D3",x"52",x"45",x"41", -- 0x0140
		x"C4",x"4C",x"45",x"D4",x"47",x"4F",x"54",x"CF", -- 0x0148
		x"52",x"55",x"CE",x"49",x"C6",x"52",x"45",x"53", -- 0x0150
		x"54",x"4F",x"52",x"C5",x"47",x"4F",x"53",x"55", -- 0x0158
		x"C2",x"52",x"45",x"54",x"55",x"52",x"CE",x"52", -- 0x0160
		x"45",x"CD",x"48",x"49",x"4D",x"45",x"CD",x"47", -- 0x0168
		x"52",x"41",x"C2",x"52",x"45",x"4C",x"45",x"41", -- 0x0170
		x"53",x"C5",x"54",x"45",x"58",x"D4",x"48",x"49", -- 0x0178
		x"52",x"45",x"D3",x"53",x"48",x"4F",x"4F",x"D4", -- 0x0180
		x"45",x"58",x"50",x"4C",x"4F",x"44",x"C5",x"5A", -- 0x0188
		x"41",x"D0",x"50",x"49",x"4E",x"C7",x"53",x"4F", -- 0x0190
		x"55",x"4E",x"C4",x"4D",x"55",x"53",x"49",x"C3", -- 0x0198
		x"50",x"4C",x"41",x"D9",x"43",x"55",x"52",x"53", -- 0x01A0
		x"45",x"D4",x"43",x"55",x"52",x"4D",x"4F",x"D6", -- 0x01A8
		x"44",x"52",x"41",x"D7",x"43",x"49",x"52",x"43", -- 0x01B0
		x"4C",x"C5",x"50",x"41",x"54",x"54",x"45",x"52", -- 0x01B8
		x"CE",x"46",x"49",x"4C",x"CC",x"43",x"48",x"41", -- 0x01C0
		x"D2",x"50",x"41",x"50",x"45",x"D2",x"49",x"4E", -- 0x01C8
		x"CB",x"53",x"54",x"4F",x"D0",x"4F",x"CE",x"57", -- 0x01D0
		x"41",x"49",x"D4",x"43",x"4C",x"4F",x"41",x"C4", -- 0x01D8
		x"43",x"53",x"41",x"56",x"C5",x"44",x"45",x"C6", -- 0x01E0
		x"50",x"4F",x"4B",x"C5",x"50",x"52",x"49",x"4E", -- 0x01E8
		x"D4",x"43",x"4F",x"4E",x"D4",x"4C",x"49",x"53", -- 0x01F0
		x"D4",x"43",x"4C",x"45",x"41",x"D2",x"47",x"45", -- 0x01F8
		x"D4",x"43",x"41",x"4C",x"CC",x"A1",x"4E",x"45", -- 0x0200
		x"D7",x"54",x"41",x"42",x"A8",x"54",x"CF",x"46", -- 0x0208
		x"CE",x"53",x"50",x"43",x"A8",x"C0",x"41",x"55", -- 0x0210
		x"54",x"CF",x"45",x"4C",x"53",x"C5",x"54",x"48", -- 0x0218
		x"45",x"CE",x"4E",x"4F",x"D4",x"53",x"54",x"45", -- 0x0220
		x"D0",x"AB",x"AD",x"AA",x"AF",x"DE",x"41",x"4E", -- 0x0228
		x"C4",x"4F",x"D2",x"BE",x"BD",x"BC",x"53",x"47", -- 0x0230
		x"CE",x"49",x"4E",x"D4",x"41",x"42",x"D3",x"55", -- 0x0238
		x"53",x"D2",x"46",x"52",x"C5",x"50",x"4F",x"D3", -- 0x0240
		x"48",x"45",x"58",x"A4",x"A6",x"53",x"51",x"D2", -- 0x0248
		x"52",x"4E",x"C4",x"4C",x"CE",x"45",x"58",x"D0", -- 0x0250
		x"43",x"4F",x"D3",x"53",x"49",x"CE",x"54",x"41", -- 0x0258
		x"CE",x"41",x"54",x"CE",x"50",x"45",x"45",x"CB", -- 0x0260
		x"44",x"45",x"45",x"CB",x"4C",x"4F",x"C7",x"4C", -- 0x0268
		x"45",x"CE",x"53",x"54",x"52",x"A4",x"56",x"41", -- 0x0270
		x"CC",x"41",x"53",x"C3",x"43",x"48",x"52",x"A4", -- 0x0278
		x"50",x"C9",x"54",x"52",x"55",x"C5",x"46",x"41", -- 0x0280
		x"4C",x"53",x"C5",x"4B",x"45",x"59",x"A4",x"53", -- 0x0288
		x"43",x"52",x"CE",x"50",x"4F",x"49",x"4E",x"D4", -- 0x0290
		x"4C",x"45",x"46",x"54",x"A4",x"52",x"49",x"47", -- 0x0298
		x"48",x"54",x"A4",x"4D",x"49",x"44",x"A4",x"00", -- 0x02A0
		x"4E",x"45",x"58",x"54",x"20",x"57",x"49",x"54", -- 0x02A8
		x"48",x"4F",x"55",x"54",x"20",x"46",x"4F",x"D2", -- 0x02B0
		x"53",x"59",x"4E",x"54",x"41",x"D8",x"52",x"45", -- 0x02B8
		x"54",x"55",x"52",x"4E",x"20",x"57",x"49",x"54", -- 0x02C0
		x"48",x"4F",x"55",x"54",x"20",x"47",x"4F",x"53", -- 0x02C8
		x"55",x"C2",x"4F",x"55",x"54",x"20",x"4F",x"46", -- 0x02D0
		x"20",x"44",x"41",x"54",x"C1",x"49",x"4C",x"4C", -- 0x02D8
		x"45",x"47",x"41",x"4C",x"20",x"51",x"55",x"41", -- 0x02E0
		x"4E",x"54",x"49",x"54",x"D9",x"4F",x"56",x"45", -- 0x02E8
		x"52",x"46",x"4C",x"4F",x"D7",x"4F",x"55",x"54", -- 0x02F0
		x"20",x"4F",x"46",x"20",x"4D",x"45",x"4D",x"4F", -- 0x02F8
		x"52",x"D9",x"55",x"4E",x"44",x"45",x"46",x"27", -- 0x0300
		x"44",x"20",x"53",x"54",x"41",x"54",x"45",x"4D", -- 0x0308
		x"45",x"4E",x"D4",x"42",x"41",x"44",x"20",x"53", -- 0x0310
		x"55",x"42",x"53",x"43",x"52",x"49",x"50",x"D4", -- 0x0318
		x"52",x"45",x"44",x"49",x"4D",x"27",x"44",x"20", -- 0x0320
		x"41",x"52",x"52",x"41",x"D9",x"44",x"49",x"56", -- 0x0328
		x"49",x"53",x"49",x"4F",x"4E",x"20",x"42",x"59", -- 0x0330
		x"20",x"5A",x"45",x"52",x"CF",x"49",x"4C",x"4C", -- 0x0338
		x"45",x"47",x"41",x"4C",x"20",x"44",x"49",x"52", -- 0x0340
		x"45",x"43",x"D4",x"44",x"49",x"53",x"50",x"20", -- 0x0348
		x"54",x"59",x"50",x"45",x"20",x"4D",x"49",x"53", -- 0x0350
		x"4D",x"41",x"54",x"43",x"C8",x"53",x"54",x"52", -- 0x0358
		x"49",x"4E",x"47",x"20",x"54",x"4F",x"4F",x"20", -- 0x0360
		x"4C",x"4F",x"4E",x"C7",x"46",x"4F",x"52",x"4D", -- 0x0368
		x"55",x"4C",x"41",x"20",x"54",x"4F",x"4F",x"20", -- 0x0370
		x"43",x"4F",x"4D",x"50",x"4C",x"45",x"D8",x"43", -- 0x0378
		x"41",x"4E",x"27",x"54",x"20",x"43",x"4F",x"4E", -- 0x0380
		x"54",x"49",x"4E",x"55",x"C5",x"55",x"4E",x"44", -- 0x0388
		x"45",x"46",x"27",x"44",x"20",x"46",x"55",x"4E", -- 0x0390
		x"43",x"54",x"49",x"4F",x"CE",x"42",x"41",x"44", -- 0x0398
		x"20",x"55",x"4E",x"54",x"49",x"CC",x"20",x"45", -- 0x03A0
		x"52",x"52",x"4F",x"52",x"00",x"20",x"49",x"4E", -- 0x03A8
		x"20",x"00",x"0D",x"0A",x"52",x"65",x"61",x"64", -- 0x03B0
		x"79",x"20",x"0D",x"0A",x"00",x"0D",x"0A",x"20", -- 0x03B8
		x"42",x"52",x"45",x"41",x"4B",x"00",x"BA",x"E8", -- 0x03C0
		x"E8",x"E8",x"E8",x"BD",x"01",x"01",x"C9",x"8D", -- 0x03C8
		x"D0",x"21",x"A5",x"B9",x"D0",x"0A",x"BD",x"02", -- 0x03D0
		x"01",x"85",x"B8",x"BD",x"03",x"01",x"85",x"B9", -- 0x03D8
		x"DD",x"03",x"01",x"D0",x"07",x"A5",x"B8",x"DD", -- 0x03E0
		x"02",x"01",x"F0",x"07",x"8A",x"18",x"69",x"12", -- 0x03E8
		x"AA",x"D0",x"D8",x"60",x"20",x"44",x"C4",x"85", -- 0x03F0
		x"A0",x"84",x"A1",x"38",x"A5",x"C9",x"E5",x"CE", -- 0x03F8
		x"85",x"91",x"A8",x"A5",x"CA",x"E5",x"CF",x"AA", -- 0x0400
		x"E8",x"98",x"F0",x"23",x"A5",x"C9",x"38",x"E5", -- 0x0408
		x"91",x"85",x"C9",x"B0",x"03",x"C6",x"CA",x"38", -- 0x0410
		x"A5",x"C7",x"E5",x"91",x"85",x"C7",x"B0",x"08", -- 0x0418
		x"C6",x"C8",x"90",x"04",x"B1",x"C9",x"91",x"C7", -- 0x0420
		x"88",x"D0",x"F9",x"B1",x"C9",x"91",x"C7",x"C6", -- 0x0428
		x"CA",x"C6",x"C8",x"CA",x"D0",x"F2",x"60",x"0A", -- 0x0430
		x"69",x"3E",x"B0",x"40",x"85",x"91",x"BA",x"E4", -- 0x0438
		x"91",x"90",x"39",x"60",x"C4",x"A3",x"90",x"28", -- 0x0440
		x"D0",x"04",x"C5",x"A2",x"90",x"22",x"48",x"A2", -- 0x0448
		x"09",x"98",x"48",x"B5",x"C6",x"CA",x"10",x"FA", -- 0x0450
		x"20",x"50",x"D6",x"A2",x"F7",x"68",x"95",x"D0", -- 0x0458
		x"E8",x"30",x"FA",x"68",x"A8",x"68",x"C4",x"A3", -- 0x0460
		x"90",x"06",x"D0",x"10",x"C5",x"A2",x"B0",x"0C", -- 0x0468
		x"60",x"AD",x"C0",x"02",x"29",x"FE",x"8D",x"C0", -- 0x0470
		x"02",x"4C",x"A8",x"C4",x"A2",x"4D",x"20",x"2F", -- 0x0478
		x"C8",x"46",x"2E",x"20",x"F0",x"CB",x"20",x"D7", -- 0x0480
		x"CC",x"BD",x"A8",x"C2",x"48",x"29",x"7F",x"20", -- 0x0488
		x"D9",x"CC",x"E8",x"68",x"10",x"F3",x"20",x"26", -- 0x0490
		x"C7",x"A9",x"A6",x"A0",x"C3",x"20",x"B0",x"CC", -- 0x0498
		x"A4",x"A9",x"C8",x"F0",x"03",x"20",x"BA",x"E0", -- 0x04A0
		x"4E",x"52",x"02",x"46",x"2E",x"4E",x"F2",x"02", -- 0x04A8
		x"A9",x"B2",x"A0",x"C3",x"20",x"1A",x"00",x"20", -- 0x04B0
		x"2F",x"C8",x"20",x"92",x"C5",x"86",x"E9",x"84", -- 0x04B8
		x"EA",x"20",x"E2",x"00",x"AA",x"F0",x"F0",x"A2", -- 0x04C0
		x"FF",x"86",x"A9",x"90",x"06",x"20",x"FA",x"C5", -- 0x04C8
		x"4C",x"0C",x"C9",x"20",x"E2",x"CA",x"20",x"FA", -- 0x04D0
		x"C5",x"84",x"26",x"20",x"B3",x"C6",x"90",x"44", -- 0x04D8
		x"A0",x"01",x"B1",x"CE",x"85",x"92",x"A5",x"9C", -- 0x04E0
		x"85",x"91",x"A5",x"CF",x"85",x"94",x"A5",x"CE", -- 0x04E8
		x"88",x"F1",x"CE",x"18",x"65",x"9C",x"85",x"9C", -- 0x04F0
		x"85",x"93",x"A5",x"9D",x"69",x"FF",x"85",x"9D", -- 0x04F8
		x"E5",x"CF",x"AA",x"38",x"A5",x"CE",x"E5",x"9C", -- 0x0500
		x"A8",x"B0",x"03",x"E8",x"C6",x"94",x"18",x"65", -- 0x0508
		x"91",x"90",x"03",x"C6",x"92",x"18",x"B1",x"91", -- 0x0510
		x"91",x"93",x"C8",x"D0",x"F9",x"E6",x"92",x"E6", -- 0x0518
		x"94",x"CA",x"D0",x"F2",x"20",x"08",x"C7",x"20", -- 0x0520
		x"5F",x"C5",x"A5",x"35",x"F0",x"89",x"18",x"A5", -- 0x0528
		x"9C",x"85",x"C9",x"65",x"26",x"85",x"C7",x"A4", -- 0x0530
		x"9D",x"84",x"CA",x"90",x"01",x"C8",x"84",x"C8", -- 0x0538
		x"20",x"F4",x"C3",x"A5",x"A0",x"A4",x"A1",x"85", -- 0x0540
		x"9C",x"84",x"9D",x"A4",x"26",x"88",x"B9",x"31", -- 0x0548
		x"00",x"91",x"CE",x"88",x"10",x"F8",x"20",x"08", -- 0x0550
		x"C7",x"20",x"5F",x"C5",x"4C",x"B7",x"C4",x"A5", -- 0x0558
		x"9A",x"A4",x"9B",x"85",x"91",x"84",x"92",x"18", -- 0x0560
		x"A0",x"01",x"B1",x"91",x"F0",x"1D",x"A0",x"04", -- 0x0568
		x"C8",x"B1",x"91",x"D0",x"FB",x"C8",x"98",x"65", -- 0x0570
		x"91",x"AA",x"A0",x"00",x"91",x"91",x"A5",x"92", -- 0x0578
		x"69",x"00",x"C8",x"91",x"91",x"86",x"91",x"85", -- 0x0580
		x"92",x"90",x"DD",x"60",x"CA",x"10",x"05",x"20", -- 0x0588
		x"F0",x"CB",x"A2",x"00",x"20",x"E8",x"C5",x"C9", -- 0x0590
		x"01",x"D0",x"0D",x"AC",x"69",x"02",x"B1",x"12", -- 0x0598
		x"29",x"7F",x"C9",x"20",x"B0",x"02",x"A9",x"09", -- 0x05A0
		x"48",x"20",x"D9",x"CC",x"68",x"C9",x"7F",x"F0", -- 0x05A8
		x"DB",x"C9",x"0D",x"F0",x"30",x"C9",x"03",x"F0", -- 0x05B0
		x"28",x"C9",x"18",x"F0",x"0B",x"C9",x"20",x"90", -- 0x05B8
		x"D3",x"95",x"35",x"E8",x"E0",x"4F",x"90",x"07", -- 0x05C0
		x"A9",x"5C",x"20",x"D9",x"CC",x"D0",x"C0",x"E0", -- 0x05C8
		x"4C",x"90",x"C1",x"8A",x"48",x"98",x"48",x"20", -- 0x05D0
		x"9F",x"FA",x"68",x"A8",x"68",x"AA",x"4C",x"94", -- 0x05D8
		x"C5",x"E6",x"17",x"A2",x"00",x"4C",x"EA",x"CB", -- 0x05E0
		x"20",x"3B",x"02",x"10",x"FB",x"C9",x"0F",x"D0", -- 0x05E8
		x"08",x"48",x"A5",x"2E",x"49",x"FF",x"85",x"2E", -- 0x05F0
		x"68",x"60",x"A6",x"E9",x"A0",x"04",x"84",x"2A", -- 0x05F8
		x"B5",x"00",x"C9",x"20",x"F0",x"41",x"85",x"25", -- 0x0600
		x"C9",x"22",x"F0",x"5F",x"24",x"2A",x"70",x"37", -- 0x0608
		x"C9",x"3F",x"D0",x"04",x"A9",x"BA",x"D0",x"2F", -- 0x0610
		x"C9",x"30",x"90",x"04",x"C9",x"3C",x"90",x"27", -- 0x0618
		x"84",x"E0",x"A0",x"00",x"84",x"26",x"A9",x"E9", -- 0x0620
		x"85",x"18",x"A9",x"C0",x"85",x"19",x"86",x"E9", -- 0x0628
		x"CA",x"E8",x"E6",x"18",x"D0",x"02",x"E6",x"19", -- 0x0630
		x"B5",x"00",x"38",x"F1",x"18",x"F0",x"F2",x"C9", -- 0x0638
		x"80",x"D0",x"2F",x"05",x"26",x"A4",x"E0",x"E8", -- 0x0640
		x"C8",x"99",x"30",x"00",x"B9",x"30",x"00",x"F0", -- 0x0648
		x"39",x"38",x"E9",x"3A",x"F0",x"04",x"C9",x"57", -- 0x0650
		x"D0",x"02",x"85",x"2A",x"38",x"E9",x"63",x"D0", -- 0x0658
		x"9F",x"85",x"25",x"B5",x"00",x"F0",x"E0",x"C5", -- 0x0660
		x"25",x"F0",x"DC",x"C8",x"99",x"30",x"00",x"E8", -- 0x0668
		x"D0",x"F1",x"A6",x"E9",x"E6",x"26",x"B1",x"18", -- 0x0670
		x"08",x"E6",x"18",x"D0",x"02",x"E6",x"19",x"28", -- 0x0678
		x"10",x"F4",x"B1",x"18",x"D0",x"B2",x"B5",x"00", -- 0x0680
		x"10",x"BB",x"99",x"32",x"00",x"A9",x"34",x"85", -- 0x0688
		x"E9",x"60",x"20",x"E2",x"CA",x"20",x"B3",x"C6", -- 0x0690
		x"90",x"16",x"6E",x"F2",x"02",x"20",x"6C",x"C7", -- 0x0698
		x"4E",x"F2",x"02",x"20",x"F0",x"CB",x"A9",x"0B", -- 0x06A0
		x"20",x"D9",x"CC",x"68",x"68",x"4C",x"B7",x"C4", -- 0x06A8
		x"4C",x"23",x"CA",x"A9",x"00",x"85",x"1D",x"85", -- 0x06B0
		x"1E",x"A5",x"9A",x"A6",x"9B",x"A0",x"01",x"85", -- 0x06B8
		x"CE",x"86",x"CF",x"B1",x"CE",x"F0",x"25",x"C8", -- 0x06C0
		x"C8",x"E6",x"1D",x"D0",x"02",x"E6",x"1E",x"A5", -- 0x06C8
		x"34",x"D1",x"CE",x"90",x"18",x"F0",x"03",x"88", -- 0x06D0
		x"D0",x"09",x"A5",x"33",x"88",x"D1",x"CE",x"90", -- 0x06D8
		x"0C",x"F0",x"0A",x"88",x"B1",x"CE",x"AA",x"88", -- 0x06E0
		x"B1",x"CE",x"B0",x"D1",x"18",x"60",x"D0",x"FD", -- 0x06E8
		x"A9",x"00",x"4E",x"F4",x"02",x"A8",x"91",x"9A", -- 0x06F0
		x"C8",x"91",x"9A",x"A5",x"9A",x"18",x"69",x"02", -- 0x06F8
		x"85",x"9C",x"A5",x"9B",x"69",x"00",x"85",x"9D", -- 0x0700
		x"20",x"3A",x"C7",x"A9",x"00",x"D0",x"2A",x"A5", -- 0x0708
		x"A6",x"A4",x"A7",x"85",x"A2",x"84",x"A3",x"A5", -- 0x0710
		x"9C",x"A4",x"9D",x"85",x"9E",x"84",x"9F",x"85", -- 0x0718
		x"A0",x"84",x"A1",x"20",x"52",x"C9",x"A2",x"88", -- 0x0720
		x"86",x"85",x"68",x"A8",x"68",x"A2",x"FE",x"9A", -- 0x0728
		x"48",x"98",x"48",x"A9",x"00",x"85",x"AD",x"85", -- 0x0730
		x"2B",x"60",x"18",x"A5",x"9A",x"69",x"FF",x"85", -- 0x0738
		x"E9",x"A5",x"9B",x"69",x"FF",x"85",x"EA",x"60", -- 0x0740
		x"08",x"20",x"E2",x"CA",x"20",x"B3",x"C6",x"28", -- 0x0748
		x"F0",x"14",x"20",x"E8",x"00",x"F0",x"15",x"C9", -- 0x0750
		x"CD",x"D0",x"92",x"20",x"E2",x"00",x"F0",x"06", -- 0x0758
		x"20",x"E2",x"CA",x"F0",x"07",x"60",x"A9",x"FF", -- 0x0760
		x"85",x"33",x"85",x"34",x"A0",x"01",x"B1",x"CE", -- 0x0768
		x"F0",x"4D",x"20",x"62",x"C9",x"C9",x"20",x"D0", -- 0x0770
		x"0E",x"4E",x"DF",x"02",x"AD",x"DF",x"02",x"10", -- 0x0778
		x"FB",x"20",x"62",x"C9",x"4E",x"DF",x"02",x"C8", -- 0x0780
		x"B1",x"CE",x"AA",x"C8",x"B1",x"CE",x"C5",x"34", -- 0x0788
		x"D0",x"04",x"E4",x"33",x"F0",x"02",x"B0",x"27", -- 0x0790
		x"84",x"B8",x"48",x"20",x"F0",x"CB",x"68",x"20", -- 0x0798
		x"C5",x"E0",x"A9",x"20",x"A4",x"B8",x"29",x"7F", -- 0x07A0
		x"20",x"D9",x"CC",x"C8",x"F0",x"11",x"B1",x"CE", -- 0x07A8
		x"D0",x"1E",x"A8",x"B1",x"CE",x"AA",x"C8",x"B1", -- 0x07B0
		x"CE",x"86",x"CE",x"85",x"CF",x"D0",x"AD",x"2C", -- 0x07B8
		x"F2",x"02",x"10",x"01",x"60",x"20",x"F0",x"CB", -- 0x07C0
		x"20",x"2F",x"C8",x"68",x"68",x"4C",x"A8",x"C4", -- 0x07C8
		x"10",x"D6",x"38",x"E9",x"7F",x"AA",x"84",x"B8", -- 0x07D0
		x"A0",x"00",x"A9",x"E9",x"85",x"18",x"A9",x"C0", -- 0x07D8
		x"85",x"19",x"CA",x"F0",x"0D",x"E6",x"18",x"D0", -- 0x07E0
		x"02",x"E6",x"19",x"B1",x"18",x"10",x"F6",x"4C", -- 0x07E8
		x"E2",x"C7",x"C8",x"B1",x"18",x"30",x"AD",x"20", -- 0x07F0
		x"D9",x"CC",x"4C",x"F2",x"C7",x"20",x"16",x"C8", -- 0x07F8
		x"4E",x"F2",x"02",x"20",x"E8",x"00",x"4C",x"48", -- 0x0800
		x"C7",x"20",x"16",x"C8",x"20",x"E8",x"00",x"20", -- 0x0808
		x"AB",x"CB",x"20",x"2F",x"C8",x"60",x"2C",x"F1", -- 0x0810
		x"02",x"30",x"39",x"A5",x"30",x"8D",x"59",x"02", -- 0x0818
		x"AD",x"58",x"02",x"85",x"30",x"38",x"6E",x"F1", -- 0x0820
		x"02",x"AD",x"56",x"02",x"4C",x"44",x"C8",x"2C", -- 0x0828
		x"F1",x"02",x"10",x"20",x"A5",x"30",x"8D",x"58", -- 0x0830
		x"02",x"AD",x"59",x"02",x"85",x"30",x"4E",x"F1", -- 0x0838
		x"02",x"AD",x"57",x"02",x"85",x"31",x"38",x"E9", -- 0x0840
		x"08",x"B0",x"FB",x"49",x"FF",x"E9",x"06",x"18", -- 0x0848
		x"65",x"31",x"85",x"32",x"60",x"A9",x"80",x"85", -- 0x0850
		x"2B",x"20",x"1C",x"CB",x"20",x"C6",x"C3",x"D0", -- 0x0858
		x"05",x"8A",x"69",x"0F",x"AA",x"9A",x"68",x"68", -- 0x0860
		x"A9",x"09",x"20",x"37",x"C4",x"20",x"4E",x"CA", -- 0x0868
		x"18",x"98",x"65",x"E9",x"48",x"A5",x"EA",x"69", -- 0x0870
		x"00",x"48",x"A5",x"A9",x"48",x"A5",x"A8",x"48", -- 0x0878
		x"A9",x"C3",x"20",x"67",x"D0",x"20",x"06",x"CF", -- 0x0880
		x"20",x"03",x"CF",x"A5",x"D5",x"09",x"7F",x"25", -- 0x0888
		x"D1",x"85",x"D1",x"A9",x"9E",x"A0",x"C8",x"85", -- 0x0890
		x"91",x"84",x"92",x"4C",x"C0",x"CF",x"A9",x"81", -- 0x0898
		x"A0",x"DC",x"20",x"7B",x"DE",x"20",x"E8",x"00", -- 0x08A0
		x"C9",x"CB",x"D0",x"06",x"20",x"E2",x"00",x"20", -- 0x08A8
		x"03",x"CF",x"20",x"13",x"DF",x"20",x"B1",x"CF", -- 0x08B0
		x"A5",x"B9",x"48",x"A5",x"B8",x"48",x"A9",x"8D", -- 0x08B8
		x"48",x"20",x"62",x"C9",x"A5",x"E9",x"A4",x"EA", -- 0x08C0
		x"F0",x"06",x"85",x"AC",x"84",x"AD",x"A0",x"00", -- 0x08C8
		x"B1",x"E9",x"D0",x"5B",x"4E",x"52",x"02",x"A0", -- 0x08D0
		x"02",x"B1",x"E9",x"18",x"D0",x"03",x"4C",x"8A", -- 0x08D8
		x"C9",x"C8",x"B1",x"E9",x"85",x"A8",x"C8",x"B1", -- 0x08E0
		x"E9",x"85",x"A9",x"98",x"65",x"E9",x"85",x"E9", -- 0x08E8
		x"90",x"02",x"E6",x"EA",x"2C",x"F4",x"02",x"10", -- 0x08F0
		x"13",x"48",x"A9",x"5B",x"20",x"FB",x"CC",x"A5", -- 0x08F8
		x"A9",x"A6",x"A8",x"20",x"C5",x"E0",x"A9",x"5D", -- 0x0900
		x"20",x"FB",x"CC",x"68",x"20",x"E2",x"00",x"20", -- 0x0908
		x"15",x"C9",x"4C",x"C1",x"C8",x"F0",x"49",x"E9", -- 0x0910
		x"80",x"90",x"11",x"C9",x"42",x"B0",x"30",x"0A", -- 0x0918
		x"A8",x"B9",x"07",x"C0",x"48",x"B9",x"06",x"C0", -- 0x0920
		x"48",x"4C",x"E2",x"00",x"4C",x"1C",x"CB",x"C9", -- 0x0928
		x"3A",x"F0",x"C1",x"C9",x"C8",x"D0",x"0E",x"2C", -- 0x0930
		x"52",x"02",x"10",x"13",x"20",x"B1",x"CA",x"4E", -- 0x0938
		x"52",x"02",x"4C",x"C1",x"C8",x"C9",x"27",x"D0", -- 0x0940
		x"06",x"20",x"99",x"CA",x"4C",x"C1",x"C8",x"4C", -- 0x0948
		x"70",x"D0",x"38",x"A5",x"9A",x"E9",x"01",x"A4", -- 0x0950
		x"9B",x"B0",x"01",x"88",x"85",x"B0",x"84",x"B1", -- 0x0958
		x"60",x"60",x"AD",x"DF",x"02",x"10",x"F9",x"29", -- 0x0960
		x"7F",x"A2",x"08",x"C9",x"03",x"D0",x"F2",x"C9", -- 0x0968
		x"03",x"B0",x"01",x"18",x"D0",x"43",x"A5",x"E9", -- 0x0970
		x"A4",x"EA",x"F0",x"0C",x"85",x"AC",x"84",x"AD", -- 0x0978
		x"A5",x"A8",x"A4",x"A9",x"85",x"AA",x"84",x"AB", -- 0x0980
		x"68",x"68",x"A9",x"BD",x"A0",x"C3",x"A2",x"00", -- 0x0988
		x"8E",x"F1",x"02",x"8E",x"DF",x"02",x"86",x"2E", -- 0x0990
		x"90",x"03",x"4C",x"9D",x"C4",x"4C",x"A8",x"C4", -- 0x0998
		x"D0",x"17",x"A2",x"D7",x"A4",x"AD",x"D0",x"03", -- 0x09A0
		x"4C",x"7E",x"C4",x"A5",x"AC",x"85",x"E9",x"84", -- 0x09A8
		x"EA",x"A5",x"AA",x"A4",x"AB",x"85",x"A8",x"84", -- 0x09B0
		x"A9",x"60",x"4C",x"36",x"D3",x"D0",x"03",x"4C", -- 0x09B8
		x"08",x"C7",x"20",x"0F",x"C7",x"4C",x"DC",x"C9", -- 0x09C0
		x"A9",x"03",x"20",x"37",x"C4",x"A5",x"EA",x"48", -- 0x09C8
		x"A5",x"E9",x"48",x"A5",x"A9",x"48",x"A5",x"A8", -- 0x09D0
		x"48",x"A9",x"9B",x"48",x"20",x"E8",x"00",x"20", -- 0x09D8
		x"E5",x"C9",x"4C",x"C1",x"C8",x"20",x"53",x"E8", -- 0x09E0
		x"20",x"51",x"CA",x"A5",x"A9",x"C5",x"34",x"B0", -- 0x09E8
		x"0B",x"98",x"38",x"65",x"E9",x"A6",x"EA",x"90", -- 0x09F0
		x"07",x"E8",x"B0",x"04",x"A5",x"9A",x"A6",x"9B", -- 0x09F8
		x"20",x"BD",x"C6",x"90",x"1E",x"A5",x"CE",x"E9", -- 0x0A00
		x"01",x"85",x"E9",x"A5",x"CF",x"E9",x"00",x"85", -- 0x0A08
		x"EA",x"60",x"D0",x"FD",x"A9",x"FF",x"85",x"B9", -- 0x0A10
		x"20",x"C6",x"C3",x"9A",x"C9",x"9B",x"F0",x"0B", -- 0x0A18
		x"A2",x"16",x"2C",x"A2",x"5A",x"4C",x"7E",x"C4", -- 0x0A20
		x"4C",x"70",x"D0",x"68",x"68",x"C0",x"0C",x"F0", -- 0x0A28
		x"19",x"85",x"A8",x"68",x"85",x"A9",x"68",x"85", -- 0x0A30
		x"E9",x"68",x"85",x"EA",x"20",x"4E",x"CA",x"98", -- 0x0A38
		x"18",x"65",x"E9",x"85",x"E9",x"90",x"02",x"E6", -- 0x0A40
		x"EA",x"60",x"68",x"68",x"68",x"60",x"A2",x"3A", -- 0x0A48
		x"2C",x"A2",x"00",x"86",x"24",x"A0",x"00",x"84", -- 0x0A50
		x"25",x"A5",x"25",x"A6",x"24",x"85",x"24",x"86", -- 0x0A58
		x"25",x"B1",x"E9",x"F0",x"E4",x"C5",x"25",x"F0", -- 0x0A60
		x"E0",x"C8",x"C9",x"22",x"D0",x"F3",x"F0",x"E9", -- 0x0A68
		x"20",x"17",x"CF",x"20",x"E8",x"00",x"C9",x"97", -- 0x0A70
		x"F0",x"05",x"A9",x"C9",x"20",x"67",x"D0",x"A5", -- 0x0A78
		x"D0",x"D0",x"05",x"20",x"9E",x"CA",x"F0",x"B7", -- 0x0A80
		x"20",x"E8",x"00",x"B0",x"03",x"4C",x"E5",x"C9", -- 0x0A88
		x"08",x"38",x"6E",x"52",x"02",x"28",x"4C",x"15", -- 0x0A90
		x"C9",x"20",x"51",x"CA",x"F0",x"A1",x"A0",x"00", -- 0x0A98
		x"B1",x"E9",x"F0",x"0C",x"C8",x"C9",x"C9",x"F0", -- 0x0AA0
		x"F0",x"C9",x"C8",x"D0",x"F3",x"4C",x"3F",x"CA", -- 0x0AA8
		x"60",x"A0",x"FF",x"C8",x"B1",x"E9",x"F0",x"04", -- 0x0AB0
		x"C9",x"3A",x"D0",x"F7",x"4C",x"3F",x"CA",x"4C", -- 0x0AB8
		x"70",x"D0",x"20",x"C8",x"D8",x"48",x"C9",x"9B", -- 0x0AC0
		x"F0",x"04",x"C9",x"97",x"D0",x"F1",x"C6",x"D4", -- 0x0AC8
		x"D0",x"04",x"68",x"4C",x"17",x"C9",x"20",x"E2", -- 0x0AD0
		x"00",x"20",x"E2",x"CA",x"C9",x"2C",x"F0",x"EE", -- 0x0AD8
		x"68",x"60",x"A2",x"00",x"86",x"33",x"86",x"34", -- 0x0AE0
		x"B0",x"F7",x"E9",x"2F",x"85",x"24",x"A5",x"34", -- 0x0AE8
		x"85",x"91",x"C9",x"19",x"B0",x"D4",x"A5",x"33", -- 0x0AF0
		x"0A",x"26",x"91",x"0A",x"26",x"91",x"65",x"33", -- 0x0AF8
		x"85",x"33",x"A5",x"91",x"65",x"34",x"85",x"34", -- 0x0B00
		x"06",x"33",x"26",x"34",x"A5",x"33",x"65",x"24", -- 0x0B08
		x"85",x"33",x"90",x"02",x"E6",x"34",x"20",x"E2", -- 0x0B10
		x"00",x"4C",x"E8",x"CA",x"20",x"88",x"D1",x"85", -- 0x0B18
		x"B8",x"84",x"B9",x"A9",x"D4",x"20",x"67",x"D0", -- 0x0B20
		x"A5",x"29",x"48",x"A5",x"28",x"48",x"20",x"17", -- 0x0B28
		x"CF",x"68",x"2A",x"20",x"09",x"CF",x"D0",x"18", -- 0x0B30
		x"68",x"10",x"12",x"20",x"F4",x"DE",x"20",x"A9", -- 0x0B38
		x"D2",x"A0",x"00",x"A5",x"D3",x"91",x"B8",x"C8", -- 0x0B40
		x"A5",x"D4",x"91",x"B8",x"60",x"4C",x"A9",x"DE", -- 0x0B48
		x"68",x"A0",x"02",x"B1",x"D3",x"C5",x"A3",x"90", -- 0x0B50
		x"17",x"D0",x"07",x"88",x"B1",x"D3",x"C5",x"A2", -- 0x0B58
		x"90",x"0E",x"A4",x"D4",x"C4",x"9D",x"90",x"08", -- 0x0B60
		x"D0",x"0D",x"A5",x"D3",x"C5",x"9C",x"B0",x"07", -- 0x0B68
		x"A5",x"D3",x"A4",x"D4",x"4C",x"8D",x"CB",x"A0", -- 0x0B70
		x"00",x"B1",x"D3",x"20",x"A3",x"D5",x"A5",x"BF", -- 0x0B78
		x"A4",x"C0",x"85",x"DE",x"84",x"DF",x"20",x"A4", -- 0x0B80
		x"D7",x"A9",x"D0",x"A0",x"00",x"85",x"BF",x"84", -- 0x0B88
		x"C0",x"20",x"05",x"D8",x"A0",x"00",x"B1",x"BF", -- 0x0B90
		x"91",x"B8",x"C8",x"B1",x"BF",x"91",x"B8",x"C8", -- 0x0B98
		x"B1",x"BF",x"91",x"B8",x"60",x"20",x"B3",x"CC", -- 0x0BA0
		x"20",x"E8",x"00",x"F0",x"43",x"F0",x"5C",x"C9", -- 0x0BA8
		x"C2",x"F0",x"7B",x"C9",x"C5",x"18",x"F0",x"76", -- 0x0BB0
		x"C9",x"2C",x"F0",x"50",x"C9",x"3B",x"F0",x"6B", -- 0x0BB8
		x"C9",x"C6",x"D0",x"03",x"4C",x"59",x"CC",x"20", -- 0x0BC0
		x"17",x"CF",x"24",x"28",x"30",x"D7",x"20",x"D5", -- 0x0BC8
		x"E0",x"20",x"B5",x"D5",x"A0",x"00",x"B1",x"D3", -- 0x0BD0
		x"18",x"65",x"30",x"C5",x"31",x"90",x"03",x"20", -- 0x0BD8
		x"F0",x"CB",x"20",x"B3",x"CC",x"20",x"D4",x"CC", -- 0x0BE0
		x"D0",x"BE",x"A0",x"00",x"94",x"35",x"A2",x"34", -- 0x0BE8
		x"A5",x"30",x"48",x"A9",x"0D",x"20",x"D9",x"CC", -- 0x0BF0
		x"68",x"2C",x"F1",x"02",x"30",x"04",x"C5",x"31", -- 0x0BF8
		x"F0",x"09",x"A9",x"00",x"85",x"30",x"A9",x"0A", -- 0x0C00
		x"20",x"D9",x"CC",x"60",x"A5",x"30",x"2C",x"F1", -- 0x0C08
		x"02",x"30",x"04",x"38",x"ED",x"53",x"02",x"38", -- 0x0C10
		x"E9",x"08",x"B0",x"FC",x"49",x"FF",x"69",x"01", -- 0x0C18
		x"AA",x"18",x"65",x"30",x"C5",x"31",x"90",x"1F", -- 0x0C20
		x"20",x"F0",x"CB",x"4C",x"4B",x"CC",x"08",x"20", -- 0x0C28
		x"C5",x"D8",x"C9",x"29",x"D0",x"20",x"28",x"90", -- 0x0C30
		x"0E",x"8A",x"C5",x"31",x"90",x"03",x"4C",x"36", -- 0x0C38
		x"D3",x"38",x"E5",x"30",x"90",x"05",x"AA",x"E8", -- 0x0C40
		x"CA",x"D0",x"06",x"20",x"E2",x"00",x"4C",x"AD", -- 0x0C48
		x"CB",x"20",x"D4",x"CC",x"D0",x"F2",x"4C",x"70", -- 0x0C50
		x"D0",x"2C",x"F1",x"02",x"30",x"F8",x"AE",x"1F", -- 0x0C58
		x"02",x"F0",x"03",x"4C",x"F7",x"EA",x"20",x"C5", -- 0x0C60
		x"D8",x"E0",x"28",x"B0",x"40",x"86",x"0C",x"20", -- 0x0C68
		x"65",x"D0",x"20",x"C8",x"D8",x"E8",x"E0",x"1C", -- 0x0C70
		x"B0",x"33",x"AD",x"6A",x"02",x"48",x"29",x"FE", -- 0x0C78
		x"8D",x"6A",x"02",x"A9",x"00",x"20",x"01",x"F8", -- 0x0C80
		x"A5",x"0C",x"8D",x"69",x"02",x"8A",x"8D",x"68", -- 0x0C88
		x"02",x"20",x"0C",x"DA",x"A5",x"1F",x"A4",x"20", -- 0x0C90
		x"85",x"12",x"84",x"13",x"68",x"8D",x"6A",x"02", -- 0x0C98
		x"A9",x"01",x"20",x"01",x"F8",x"A9",x"3B",x"20", -- 0x0CA0
		x"67",x"D0",x"4C",x"AD",x"CB",x"4C",x"C2",x"D8", -- 0x0CA8
		x"20",x"B5",x"D5",x"20",x"D0",x"D7",x"AA",x"A0", -- 0x0CB0
		x"00",x"E8",x"CA",x"F0",x"10",x"B1",x"91",x"20", -- 0x0CB8
		x"D9",x"CC",x"C8",x"C9",x"0D",x"D0",x"F3",x"20", -- 0x0CC0
		x"0B",x"CC",x"4C",x"BA",x"CC",x"60",x"A9",x"0C", -- 0x0CC8
		x"2C",x"A9",x"11",x"2C",x"A9",x"20",x"2C",x"A9", -- 0x0CD0
		x"3F",x"24",x"2E",x"30",x"33",x"48",x"C9",x"20", -- 0x0CD8
		x"90",x"0B",x"A5",x"30",x"C5",x"31",x"D0",x"03", -- 0x0CE0
		x"20",x"F0",x"CB",x"E6",x"30",x"68",x"2C",x"F1", -- 0x0CE8
		x"02",x"10",x"08",x"48",x"20",x"3E",x"02",x"68", -- 0x0CF0
		x"29",x"FF",x"60",x"86",x"27",x"AA",x"20",x"7C", -- 0x0CF8
		x"F7",x"C9",x"20",x"90",x"04",x"C9",x"7F",x"D0", -- 0x0D00
		x"05",x"AE",x"69",x"02",x"86",x"30",x"A6",x"27", -- 0x0D08
		x"29",x"FF",x"60",x"6C",x"F5",x"02",x"A9",x"80", -- 0x0D10
		x"2C",x"A9",x"00",x"8D",x"F4",x"02",x"60",x"A5", -- 0x0D18
		x"2C",x"F0",x"13",x"30",x"04",x"A0",x"FF",x"D0", -- 0x0D20
		x"04",x"A5",x"AE",x"A4",x"AF",x"85",x"A8",x"84", -- 0x0D28
		x"A9",x"A2",x"A8",x"4C",x"7E",x"C4",x"A9",x"85", -- 0x0D30
		x"A0",x"CE",x"20",x"B0",x"CC",x"A5",x"AC",x"A4", -- 0x0D38
		x"AD",x"85",x"E9",x"84",x"EA",x"60",x"20",x"D2", -- 0x0D40
		x"D4",x"A2",x"36",x"A0",x"00",x"84",x"36",x"A9", -- 0x0D48
		x"40",x"20",x"8F",x"CD",x"60",x"46",x"2E",x"C9", -- 0x0D50
		x"22",x"D0",x"0B",x"20",x"25",x"D0",x"A9",x"3B", -- 0x0D58
		x"20",x"67",x"D0",x"20",x"B3",x"CC",x"20",x"D2", -- 0x0D60
		x"D4",x"A9",x"2C",x"85",x"34",x"A9",x"00",x"85", -- 0x0D68
		x"17",x"20",x"80",x"CD",x"A5",x"35",x"D0",x"16", -- 0x0D70
		x"A5",x"17",x"F0",x"F1",x"18",x"4C",x"80",x"C9", -- 0x0D78
		x"20",x"D7",x"CC",x"20",x"D4",x"CC",x"4C",x"92", -- 0x0D80
		x"C5",x"A6",x"B0",x"A4",x"B1",x"A9",x"98",x"85", -- 0x0D88
		x"2C",x"86",x"B2",x"84",x"B3",x"20",x"88",x"D1", -- 0x0D90
		x"85",x"B8",x"84",x"B9",x"A5",x"E9",x"A4",x"EA", -- 0x0D98
		x"85",x"BA",x"84",x"BB",x"A6",x"B2",x"A4",x"B3", -- 0x0DA0
		x"86",x"E9",x"84",x"EA",x"20",x"E8",x"00",x"D0", -- 0x0DA8
		x"1D",x"24",x"2C",x"50",x"0D",x"20",x"78",x"EB", -- 0x0DB0
		x"10",x"FB",x"85",x"35",x"A2",x"34",x"A0",x"00", -- 0x0DB8
		x"F0",x"08",x"30",x"71",x"20",x"D7",x"CC",x"20", -- 0x0DC0
		x"80",x"CD",x"86",x"E9",x"84",x"EA",x"20",x"E2", -- 0x0DC8
		x"00",x"24",x"28",x"10",x"31",x"24",x"2C",x"50", -- 0x0DD0
		x"09",x"E8",x"86",x"E9",x"A9",x"00",x"85",x"24", -- 0x0DD8
		x"F0",x"0C",x"85",x"24",x"C9",x"22",x"F0",x"07", -- 0x0DE0
		x"A9",x"3A",x"85",x"24",x"A9",x"2C",x"18",x"85", -- 0x0DE8
		x"25",x"A5",x"E9",x"A4",x"EA",x"69",x"00",x"90", -- 0x0DF0
		x"01",x"C8",x"20",x"BB",x"D5",x"20",x"0D",x"D9", -- 0x0DF8
		x"20",x"51",x"CB",x"4C",x"0E",x"CE",x"20",x"E7", -- 0x0E00
		x"DF",x"A5",x"29",x"20",x"39",x"CB",x"20",x"E8", -- 0x0E08
		x"00",x"F0",x"07",x"C9",x"2C",x"F0",x"03",x"4C", -- 0x0E10
		x"1F",x"CD",x"A5",x"E9",x"A4",x"EA",x"85",x"B2", -- 0x0E18
		x"84",x"B3",x"A5",x"BA",x"A4",x"BB",x"85",x"E9", -- 0x0E20
		x"84",x"EA",x"20",x"E8",x"00",x"F0",x"2C",x"20", -- 0x0E28
		x"65",x"D0",x"4C",x"95",x"CD",x"20",x"4E",x"CA", -- 0x0E30
		x"C8",x"AA",x"D0",x"12",x"A2",x"2A",x"C8",x"B1", -- 0x0E38
		x"E9",x"F0",x"69",x"C8",x"B1",x"E9",x"85",x"AE", -- 0x0E40
		x"C8",x"B1",x"E9",x"C8",x"85",x"AF",x"B1",x"E9", -- 0x0E48
		x"AA",x"20",x"3F",x"CA",x"E0",x"91",x"D0",x"DD", -- 0x0E50
		x"4C",x"CE",x"CD",x"A5",x"B2",x"A4",x"B3",x"A6", -- 0x0E58
		x"2C",x"10",x"03",x"4C",x"5C",x"C9",x"A0",x"00", -- 0x0E60
		x"B1",x"B2",x"F0",x"07",x"A9",x"74",x"A0",x"CE", -- 0x0E68
		x"4C",x"B0",x"CC",x"60",x"3F",x"45",x"58",x"54", -- 0x0E70
		x"52",x"41",x"20",x"49",x"47",x"4E",x"4F",x"52", -- 0x0E78
		x"45",x"44",x"0D",x"0A",x"00",x"3F",x"52",x"45", -- 0x0E80
		x"44",x"4F",x"20",x"46",x"52",x"4F",x"4D",x"20", -- 0x0E88
		x"53",x"54",x"41",x"52",x"54",x"0D",x"0A",x"00", -- 0x0E90
		x"D0",x"04",x"A0",x"00",x"F0",x"03",x"20",x"88", -- 0x0E98
		x"D1",x"85",x"B8",x"84",x"B9",x"20",x"C6",x"C3", -- 0x0EA0
		x"F0",x"04",x"A2",x"00",x"F0",x"66",x"9A",x"8A", -- 0x0EA8
		x"18",x"69",x"04",x"48",x"69",x"06",x"85",x"93", -- 0x0EB0
		x"68",x"A0",x"01",x"20",x"7B",x"DE",x"BA",x"BD", -- 0x0EB8
		x"09",x"01",x"85",x"D5",x"A5",x"B8",x"A4",x"B9", -- 0x0EC0
		x"20",x"22",x"DB",x"20",x"A9",x"DE",x"A0",x"01", -- 0x0EC8
		x"20",x"4E",x"DF",x"BA",x"38",x"FD",x"09",x"01", -- 0x0ED0
		x"F0",x"17",x"BD",x"0F",x"01",x"85",x"A8",x"BD", -- 0x0ED8
		x"10",x"01",x"85",x"A9",x"BD",x"12",x"01",x"85", -- 0x0EE0
		x"E9",x"BD",x"11",x"01",x"85",x"EA",x"4C",x"C1", -- 0x0EE8
		x"C8",x"8A",x"69",x"11",x"AA",x"9A",x"20",x"E8", -- 0x0EF0
		x"00",x"C9",x"2C",x"D0",x"F1",x"20",x"E2",x"00", -- 0x0EF8
		x"20",x"9E",x"CE",x"20",x"17",x"CF",x"18",x"24", -- 0x0F00
		x"38",x"24",x"28",x"30",x"03",x"B0",x"03",x"60", -- 0x0F08
		x"B0",x"FD",x"A2",x"A8",x"4C",x"7E",x"C4",x"A6", -- 0x0F10
		x"E9",x"D0",x"02",x"C6",x"EA",x"C6",x"E9",x"A2", -- 0x0F18
		x"00",x"24",x"48",x"8A",x"48",x"A9",x"01",x"20", -- 0x0F20
		x"37",x"C4",x"20",x"00",x"D0",x"A9",x"00",x"85", -- 0x0F28
		x"BC",x"20",x"E8",x"00",x"38",x"E9",x"D3",x"90", -- 0x0F30
		x"17",x"C9",x"03",x"B0",x"13",x"C9",x"01",x"2A", -- 0x0F38
		x"49",x"01",x"45",x"BC",x"C5",x"BC",x"90",x"61", -- 0x0F40
		x"85",x"BC",x"20",x"E2",x"00",x"4C",x"34",x"CF", -- 0x0F48
		x"A6",x"BC",x"D0",x"2C",x"B0",x"7F",x"69",x"07", -- 0x0F50
		x"90",x"7B",x"65",x"28",x"D0",x"03",x"4C",x"67", -- 0x0F58
		x"D7",x"69",x"FF",x"85",x"91",x"0A",x"65",x"91", -- 0x0F60
		x"A8",x"68",x"D9",x"CC",x"C0",x"B0",x"6B",x"20", -- 0x0F68
		x"06",x"CF",x"48",x"20",x"99",x"CF",x"68",x"A4", -- 0x0F70
		x"BA",x"10",x"17",x"AA",x"F0",x"5A",x"D0",x"63", -- 0x0F78
		x"46",x"28",x"8A",x"2A",x"A6",x"E9",x"D0",x"02", -- 0x0F80
		x"C6",x"EA",x"C6",x"E9",x"A0",x"1B",x"85",x"BC", -- 0x0F88
		x"D0",x"D7",x"D9",x"CC",x"C0",x"B0",x"4C",x"90", -- 0x0F90
		x"D9",x"B9",x"CE",x"C0",x"48",x"B9",x"CD",x"C0", -- 0x0F98
		x"48",x"20",x"AC",x"CF",x"A5",x"BC",x"4C",x"22", -- 0x0FA0
		x"CF",x"4C",x"70",x"D0",x"A5",x"D5",x"BE",x"CC", -- 0x0FA8
		x"C0",x"A8",x"68",x"85",x"91",x"68",x"85",x"92", -- 0x0FB0
		x"E6",x"91",x"D0",x"02",x"E6",x"92",x"98",x"48", -- 0x0FB8
		x"20",x"F4",x"DE",x"A5",x"D4",x"48",x"A5",x"D3", -- 0x0FC0
		x"48",x"A5",x"D2",x"48",x"A5",x"D1",x"48",x"A5", -- 0x0FC8
		x"D0",x"48",x"6C",x"91",x"00",x"A0",x"FF",x"68", -- 0x0FD0
		x"F0",x"23",x"C9",x"64",x"F0",x"03",x"20",x"06", -- 0x0FD8
		x"CF",x"84",x"BA",x"68",x"4A",x"85",x"2D",x"68", -- 0x0FE0
		x"85",x"D8",x"68",x"85",x"D9",x"68",x"85",x"DA", -- 0x0FE8
		x"68",x"85",x"DB",x"68",x"85",x"DC",x"68",x"85", -- 0x0FF0
		x"DD",x"45",x"D5",x"85",x"DE",x"A5",x"D0",x"60", -- 0x0FF8
		x"A9",x"00",x"85",x"28",x"20",x"E2",x"00",x"B0", -- 0x1000
		x"03",x"4C",x"E7",x"DF",x"20",x"16",x"D2",x"B0", -- 0x1008
		x"6B",x"C9",x"2E",x"F0",x"F4",x"C9",x"23",x"F0", -- 0x1010
		x"F0",x"C9",x"CD",x"F0",x"58",x"C9",x"CC",x"F0", -- 0x1018
		x"E3",x"C9",x"22",x"D0",x"0F",x"A5",x"E9",x"A4", -- 0x1020
		x"EA",x"69",x"00",x"90",x"01",x"C8",x"20",x"B5", -- 0x1028
		x"D5",x"4C",x"0D",x"D9",x"C9",x"CA",x"D0",x"13", -- 0x1030
		x"A0",x"18",x"D0",x"3B",x"20",x"A9",x"D2",x"A5", -- 0x1038
		x"D4",x"49",x"FF",x"A8",x"A5",x"D3",x"49",x"FF", -- 0x1040
		x"4C",x"99",x"D4",x"C9",x"C4",x"D0",x"03",x"4C", -- 0x1048
		x"22",x"D5",x"C9",x"D6",x"90",x"03",x"4C",x"A0", -- 0x1050
		x"D0",x"20",x"62",x"D0",x"20",x"17",x"CF",x"A9", -- 0x1058
		x"29",x"2C",x"A9",x"28",x"2C",x"A9",x"2C",x"A0", -- 0x1060
		x"00",x"D1",x"E9",x"D0",x"03",x"4C",x"E2",x"00", -- 0x1068
		x"A2",x"10",x"4C",x"7E",x"C4",x"A0",x"15",x"68", -- 0x1070
		x"68",x"4C",x"73",x"CF",x"20",x"88",x"D1",x"85", -- 0x1078
		x"D3",x"84",x"D4",x"A6",x"28",x"F0",x"05",x"A2", -- 0x1080
		x"00",x"86",x"DF",x"60",x"A6",x"29",x"10",x"0D", -- 0x1088
		x"A0",x"00",x"B1",x"D3",x"AA",x"C8",x"B1",x"D3", -- 0x1090
		x"A8",x"8A",x"4C",x"99",x"D4",x"4C",x"7B",x"DE", -- 0x1098
		x"0A",x"48",x"AA",x"20",x"E2",x"00",x"E0",x"DB", -- 0x10A0
		x"90",x"24",x"E0",x"E7",x"90",x"23",x"20",x"62", -- 0x10A8
		x"D0",x"20",x"17",x"CF",x"20",x"65",x"D0",x"20", -- 0x10B0
		x"08",x"CF",x"68",x"AA",x"A5",x"D4",x"48",x"A5", -- 0x10B8
		x"D3",x"48",x"8A",x"48",x"20",x"C8",x"D8",x"68", -- 0x10C0
		x"A8",x"8A",x"48",x"4C",x"D3",x"D0",x"20",x"59", -- 0x10C8
		x"D0",x"68",x"A8",x"B9",x"DE",x"BF",x"85",x"C4", -- 0x10D0
		x"B9",x"DF",x"BF",x"85",x"C5",x"20",x"C3",x"00", -- 0x10D8
		x"4C",x"06",x"CF",x"A0",x"FF",x"2C",x"A0",x"00", -- 0x10E0
		x"84",x"26",x"20",x"A9",x"D2",x"A5",x"D3",x"45", -- 0x10E8
		x"26",x"85",x"24",x"A5",x"D4",x"45",x"26",x"85", -- 0x10F0
		x"25",x"20",x"D5",x"DE",x"20",x"A9",x"D2",x"A5", -- 0x10F8
		x"D4",x"45",x"26",x"25",x"25",x"45",x"26",x"A8", -- 0x1100
		x"A5",x"D3",x"45",x"26",x"25",x"24",x"45",x"26", -- 0x1108
		x"4C",x"99",x"D4",x"20",x"09",x"CF",x"B0",x"13", -- 0x1110
		x"A5",x"DD",x"09",x"7F",x"25",x"D9",x"85",x"D9", -- 0x1118
		x"A9",x"D8",x"A0",x"00",x"20",x"4C",x"DF",x"AA", -- 0x1120
		x"4C",x"5E",x"D1",x"A9",x"00",x"85",x"28",x"C6", -- 0x1128
		x"BC",x"20",x"D0",x"D7",x"85",x"D0",x"86",x"D1", -- 0x1130
		x"84",x"D2",x"A5",x"DB",x"A4",x"DC",x"20",x"D4", -- 0x1138
		x"D7",x"86",x"DB",x"84",x"DC",x"AA",x"38",x"E5", -- 0x1140
		x"D0",x"F0",x"08",x"A9",x"01",x"90",x"04",x"A6", -- 0x1148
		x"D0",x"A9",x"FF",x"85",x"D5",x"A0",x"FF",x"E8", -- 0x1150
		x"C8",x"CA",x"D0",x"07",x"A6",x"D5",x"30",x"0F", -- 0x1158
		x"18",x"90",x"0C",x"B1",x"DB",x"D1",x"D1",x"F0", -- 0x1160
		x"EF",x"A2",x"FF",x"B0",x"02",x"A2",x"01",x"E8", -- 0x1168
		x"8A",x"2A",x"25",x"2D",x"F0",x"02",x"A9",x"FF", -- 0x1170
		x"4C",x"24",x"DF",x"20",x"65",x"D0",x"AA",x"20", -- 0x1178
		x"8D",x"D1",x"20",x"E8",x"00",x"D0",x"F4",x"60", -- 0x1180
		x"A2",x"00",x"20",x"E8",x"00",x"86",x"27",x"85", -- 0x1188
		x"B4",x"20",x"E8",x"00",x"20",x"16",x"D2",x"B0", -- 0x1190
		x"03",x"4C",x"70",x"D0",x"A2",x"00",x"86",x"28", -- 0x1198
		x"86",x"29",x"20",x"E2",x"00",x"90",x"05",x"20", -- 0x11A0
		x"16",x"D2",x"90",x"0B",x"AA",x"20",x"E2",x"00", -- 0x11A8
		x"90",x"FB",x"20",x"16",x"D2",x"B0",x"F6",x"C9", -- 0x11B0
		x"24",x"D0",x"06",x"A9",x"FF",x"85",x"28",x"D0", -- 0x11B8
		x"10",x"C9",x"25",x"D0",x"13",x"A5",x"2B",x"30", -- 0x11C0
		x"D0",x"A9",x"80",x"85",x"29",x"05",x"B4",x"85", -- 0x11C8
		x"B4",x"8A",x"09",x"80",x"AA",x"20",x"E2",x"00", -- 0x11D0
		x"86",x"B5",x"38",x"05",x"2B",x"E9",x"28",x"D0", -- 0x11D8
		x"03",x"4C",x"BB",x"D2",x"24",x"2B",x"70",x"F9", -- 0x11E0
		x"A9",x"00",x"85",x"2B",x"A5",x"9C",x"A6",x"9D", -- 0x11E8
		x"A0",x"00",x"86",x"CF",x"85",x"CE",x"E4",x"9F", -- 0x11F0
		x"D0",x"04",x"C5",x"9E",x"F0",x"24",x"A5",x"B4", -- 0x11F8
		x"D1",x"CE",x"D0",x"08",x"A5",x"B5",x"C8",x"D1", -- 0x1200
		x"CE",x"F0",x"6C",x"88",x"18",x"A5",x"CE",x"69", -- 0x1208
		x"07",x"90",x"E1",x"E8",x"D0",x"DC",x"C9",x"41", -- 0x1210
		x"90",x"07",x"E9",x"5B",x"38",x"E9",x"A5",x"B0", -- 0x1218
		x"00",x"60",x"68",x"48",x"C9",x"7E",x"D0",x"0D", -- 0x1220
		x"BA",x"BD",x"02",x"01",x"C9",x"D0",x"D0",x"05", -- 0x1228
		x"A9",x"07",x"A0",x"E2",x"60",x"A5",x"9E",x"A4", -- 0x1230
		x"9F",x"85",x"CE",x"84",x"CF",x"A5",x"A0",x"A4", -- 0x1238
		x"A1",x"85",x"C9",x"84",x"CA",x"18",x"69",x"07", -- 0x1240
		x"90",x"01",x"C8",x"85",x"C7",x"84",x"C8",x"20", -- 0x1248
		x"F4",x"C3",x"A5",x"C7",x"A4",x"C8",x"C8",x"85", -- 0x1250
		x"9E",x"84",x"9F",x"A0",x"00",x"A5",x"B4",x"91", -- 0x1258
		x"CE",x"C8",x"A5",x"B5",x"91",x"CE",x"A9",x"00", -- 0x1260
		x"C8",x"91",x"CE",x"C8",x"91",x"CE",x"C8",x"91", -- 0x1268
		x"CE",x"C8",x"91",x"CE",x"C8",x"91",x"CE",x"A5", -- 0x1270
		x"CE",x"18",x"69",x"02",x"A4",x"CF",x"90",x"01", -- 0x1278
		x"C8",x"85",x"B6",x"84",x"B7",x"60",x"A5",x"26", -- 0x1280
		x"0A",x"69",x"05",x"65",x"CE",x"A4",x"CF",x"90", -- 0x1288
		x"01",x"C8",x"85",x"C7",x"84",x"C8",x"60",x"90", -- 0x1290
		x"80",x"00",x"00",x"00",x"20",x"E2",x"00",x"20", -- 0x1298
		x"17",x"CF",x"20",x"06",x"CF",x"A5",x"D5",x"30", -- 0x12A0
		x"0D",x"A5",x"D0",x"C9",x"90",x"90",x"09",x"A9", -- 0x12A8
		x"97",x"A0",x"D2",x"20",x"4C",x"DF",x"D0",x"7E", -- 0x12B0
		x"4C",x"8C",x"DF",x"A5",x"2B",x"D0",x"47",x"A5", -- 0x12B8
		x"27",x"05",x"29",x"48",x"A5",x"28",x"48",x"A0", -- 0x12C0
		x"00",x"98",x"48",x"A5",x"B5",x"48",x"A5",x"B4", -- 0x12C8
		x"48",x"20",x"9C",x"D2",x"68",x"85",x"B4",x"68", -- 0x12D0
		x"85",x"B5",x"68",x"A8",x"BA",x"BD",x"02",x"01", -- 0x12D8
		x"48",x"BD",x"01",x"01",x"48",x"A5",x"D3",x"9D", -- 0x12E0
		x"02",x"01",x"A5",x"D4",x"9D",x"01",x"01",x"C8", -- 0x12E8
		x"20",x"E8",x"00",x"C9",x"2C",x"F0",x"D2",x"84", -- 0x12F0
		x"26",x"20",x"5F",x"D0",x"68",x"85",x"28",x"68", -- 0x12F8
		x"85",x"29",x"29",x"7F",x"85",x"27",x"A6",x"9E", -- 0x1300
		x"A5",x"9F",x"86",x"CE",x"85",x"CF",x"C5",x"A1", -- 0x1308
		x"D0",x"04",x"E4",x"A0",x"F0",x"3F",x"A0",x"00", -- 0x1310
		x"B1",x"CE",x"C8",x"C5",x"B4",x"D0",x"06",x"A5", -- 0x1318
		x"B5",x"D1",x"CE",x"F0",x"16",x"C8",x"B1",x"CE", -- 0x1320
		x"18",x"65",x"CE",x"AA",x"C8",x"B1",x"CE",x"65", -- 0x1328
		x"CF",x"90",x"D7",x"A2",x"6B",x"2C",x"A2",x"35", -- 0x1330
		x"4C",x"7E",x"C4",x"A2",x"78",x"A5",x"27",x"D0", -- 0x1338
		x"F7",x"A5",x"2B",x"F0",x"02",x"38",x"60",x"20", -- 0x1340
		x"86",x"D2",x"A5",x"26",x"A0",x"04",x"D1",x"CE", -- 0x1348
		x"D0",x"E1",x"4C",x"EB",x"D3",x"A5",x"2B",x"F0", -- 0x1350
		x"08",x"20",x"3D",x"E9",x"A2",x"2A",x"4C",x"7E", -- 0x1358
		x"C4",x"20",x"86",x"D2",x"20",x"44",x"C4",x"A9", -- 0x1360
		x"00",x"A8",x"85",x"E1",x"A2",x"05",x"A5",x"B4", -- 0x1368
		x"91",x"CE",x"10",x"01",x"CA",x"C8",x"A5",x"B5", -- 0x1370
		x"91",x"CE",x"10",x"02",x"CA",x"CA",x"86",x"E0", -- 0x1378
		x"A5",x"26",x"C8",x"C8",x"C8",x"91",x"CE",x"A2", -- 0x1380
		x"0B",x"A9",x"00",x"24",x"27",x"50",x"08",x"68", -- 0x1388
		x"18",x"69",x"01",x"AA",x"68",x"69",x"00",x"C8", -- 0x1390
		x"91",x"CE",x"C8",x"8A",x"91",x"CE",x"20",x"4D", -- 0x1398
		x"D4",x"86",x"E0",x"85",x"E1",x"A4",x"91",x"C6", -- 0x13A0
		x"26",x"D0",x"DC",x"65",x"C8",x"B0",x"5D",x"85", -- 0x13A8
		x"C8",x"A8",x"8A",x"65",x"C7",x"90",x"03",x"C8", -- 0x13B0
		x"F0",x"52",x"20",x"44",x"C4",x"85",x"A0",x"84", -- 0x13B8
		x"A1",x"A9",x"00",x"E6",x"E1",x"A4",x"E0",x"F0", -- 0x13C0
		x"05",x"88",x"91",x"C7",x"D0",x"FB",x"C6",x"C8", -- 0x13C8
		x"C6",x"E1",x"D0",x"F5",x"E6",x"C8",x"38",x"A5", -- 0x13D0
		x"A0",x"E5",x"CE",x"A0",x"02",x"91",x"CE",x"A5", -- 0x13D8
		x"A1",x"C8",x"E5",x"CF",x"91",x"CE",x"A5",x"27", -- 0x13E0
		x"D0",x"62",x"C8",x"B1",x"CE",x"85",x"26",x"A9", -- 0x13E8
		x"00",x"85",x"E0",x"85",x"E1",x"C8",x"68",x"AA", -- 0x13F0
		x"85",x"D3",x"68",x"85",x"D4",x"D1",x"CE",x"90", -- 0x13F8
		x"0E",x"D0",x"06",x"C8",x"8A",x"D1",x"CE",x"90", -- 0x1400
		x"07",x"4C",x"33",x"D3",x"4C",x"7C",x"C4",x"C8", -- 0x1408
		x"A5",x"E1",x"05",x"E0",x"18",x"F0",x"0A",x"20", -- 0x1410
		x"4D",x"D4",x"8A",x"65",x"D3",x"AA",x"98",x"A4", -- 0x1418
		x"91",x"65",x"D4",x"86",x"E0",x"C6",x"26",x"D0", -- 0x1420
		x"CA",x"85",x"E1",x"A2",x"05",x"A5",x"B4",x"10", -- 0x1428
		x"01",x"CA",x"A5",x"B5",x"10",x"02",x"CA",x"CA", -- 0x1430
		x"86",x"97",x"A9",x"00",x"20",x"56",x"D4",x"8A", -- 0x1438
		x"65",x"C7",x"85",x"B6",x"98",x"65",x"C8",x"85", -- 0x1440
		x"B7",x"A8",x"A5",x"B6",x"60",x"84",x"91",x"B1", -- 0x1448
		x"CE",x"85",x"97",x"88",x"B1",x"CE",x"85",x"98", -- 0x1450
		x"A9",x"10",x"85",x"CC",x"A2",x"00",x"A0",x"00", -- 0x1458
		x"8A",x"0A",x"AA",x"98",x"2A",x"A8",x"B0",x"A4", -- 0x1460
		x"06",x"E0",x"26",x"E1",x"90",x"0B",x"18",x"8A", -- 0x1468
		x"65",x"97",x"AA",x"98",x"65",x"98",x"A8",x"B0", -- 0x1470
		x"93",x"C6",x"CC",x"D0",x"E3",x"60",x"A5",x"28", -- 0x1478
		x"F0",x"03",x"20",x"D0",x"D7",x"20",x"50",x"D6", -- 0x1480
		x"38",x"A5",x"A2",x"E5",x"A0",x"A8",x"A5",x"A3", -- 0x1488
		x"E5",x"A1",x"A2",x"00",x"86",x"28",x"4C",x"40", -- 0x1490
		x"DF",x"A2",x"00",x"86",x"28",x"85",x"D1",x"84", -- 0x1498
		x"D2",x"A2",x"90",x"4C",x"2C",x"DF",x"20",x"CB", -- 0x14A0
		x"D8",x"8A",x"F0",x"08",x"AC",x"58",x"02",x"2C", -- 0x14A8
		x"F1",x"02",x"10",x"02",x"A4",x"30",x"A9",x"00", -- 0x14B0
		x"F0",x"DF",x"C9",x"D9",x"D0",x"21",x"20",x"E2", -- 0x14B8
		x"00",x"A9",x"D4",x"20",x"67",x"D0",x"20",x"53", -- 0x14C0
		x"E8",x"A5",x"33",x"A4",x"34",x"85",x"22",x"84", -- 0x14C8
		x"23",x"60",x"A6",x"A9",x"E8",x"D0",x"FA",x"A2", -- 0x14D0
		x"95",x"2C",x"A2",x"E5",x"4C",x"7E",x"C4",x"20", -- 0x14D8
		x"0D",x"D5",x"20",x"D2",x"D4",x"20",x"62",x"D0", -- 0x14E0
		x"A9",x"80",x"85",x"2B",x"20",x"88",x"D1",x"20", -- 0x14E8
		x"06",x"CF",x"20",x"5F",x"D0",x"A9",x"D4",x"20", -- 0x14F0
		x"67",x"D0",x"48",x"A5",x"B7",x"48",x"A5",x"B6", -- 0x14F8
		x"48",x"A5",x"EA",x"48",x"A5",x"E9",x"48",x"20", -- 0x1500
		x"3C",x"CA",x"4C",x"7D",x"D5",x"A9",x"C4",x"20", -- 0x1508
		x"67",x"D0",x"09",x"80",x"A2",x"80",x"86",x"2B", -- 0x1510
		x"20",x"8F",x"D1",x"85",x"BD",x"84",x"BE",x"4C", -- 0x1518
		x"06",x"CF",x"20",x"0D",x"D5",x"A5",x"BE",x"48", -- 0x1520
		x"A5",x"BD",x"48",x"20",x"59",x"D0",x"20",x"06", -- 0x1528
		x"CF",x"68",x"85",x"BD",x"68",x"85",x"BE",x"A0", -- 0x1530
		x"02",x"B1",x"BD",x"85",x"B6",x"AA",x"C8",x"B1", -- 0x1538
		x"BD",x"F0",x"97",x"85",x"B7",x"C8",x"B1",x"B6", -- 0x1540
		x"48",x"88",x"10",x"FA",x"A4",x"B7",x"20",x"AD", -- 0x1548
		x"DE",x"A5",x"EA",x"48",x"A5",x"E9",x"48",x"B1", -- 0x1550
		x"BD",x"85",x"E9",x"C8",x"B1",x"BD",x"85",x"EA", -- 0x1558
		x"A5",x"B7",x"48",x"A5",x"B6",x"48",x"20",x"03", -- 0x1560
		x"CF",x"68",x"85",x"BD",x"68",x"85",x"BE",x"20", -- 0x1568
		x"E8",x"00",x"F0",x"03",x"4C",x"70",x"D0",x"68", -- 0x1570
		x"85",x"E9",x"68",x"85",x"EA",x"A0",x"00",x"68", -- 0x1578
		x"91",x"BD",x"68",x"C8",x"91",x"BD",x"68",x"C8", -- 0x1580
		x"91",x"BD",x"68",x"C8",x"91",x"BD",x"68",x"C8", -- 0x1588
		x"91",x"BD",x"60",x"20",x"06",x"CF",x"A0",x"00", -- 0x1590
		x"20",x"D7",x"E0",x"68",x"68",x"A9",x"FF",x"A0", -- 0x1598
		x"00",x"F0",x"12",x"A6",x"D3",x"A4",x"D4",x"86", -- 0x15A0
		x"BF",x"84",x"C0",x"20",x"1E",x"D6",x"86",x"D1", -- 0x15A8
		x"84",x"D2",x"85",x"D0",x"60",x"A2",x"22",x"86", -- 0x15B0
		x"24",x"86",x"25",x"85",x"DE",x"84",x"DF",x"85", -- 0x15B8
		x"D1",x"84",x"D2",x"A0",x"FF",x"C8",x"B1",x"DE", -- 0x15C0
		x"F0",x"0C",x"C5",x"24",x"F0",x"04",x"C5",x"25", -- 0x15C8
		x"D0",x"F3",x"C9",x"22",x"F0",x"01",x"18",x"84", -- 0x15D0
		x"D0",x"98",x"65",x"DE",x"85",x"E0",x"A6",x"DF", -- 0x15D8
		x"90",x"01",x"E8",x"86",x"E1",x"A5",x"DF",x"D0", -- 0x15E0
		x"0B",x"98",x"20",x"A3",x"D5",x"A6",x"DE",x"A4", -- 0x15E8
		x"DF",x"20",x"B2",x"D7",x"A6",x"85",x"E0",x"91", -- 0x15F0
		x"D0",x"05",x"A2",x"C4",x"4C",x"7E",x"C4",x"A5", -- 0x15F8
		x"D0",x"95",x"00",x"A5",x"D1",x"95",x"01",x"A5", -- 0x1600
		x"D2",x"95",x"02",x"A0",x"00",x"86",x"D3",x"84", -- 0x1608
		x"D4",x"84",x"DF",x"88",x"84",x"28",x"86",x"86", -- 0x1610
		x"E8",x"E8",x"E8",x"86",x"85",x"60",x"46",x"2A", -- 0x1618
		x"48",x"49",x"FF",x"38",x"65",x"A2",x"A4",x"A3", -- 0x1620
		x"B0",x"01",x"88",x"C4",x"A1",x"90",x"11",x"D0", -- 0x1628
		x"04",x"C5",x"A0",x"90",x"0B",x"85",x"A2",x"84", -- 0x1630
		x"A3",x"85",x"A4",x"84",x"A5",x"AA",x"68",x"60", -- 0x1638
		x"A2",x"4D",x"A5",x"2A",x"30",x"B6",x"20",x"50", -- 0x1640
		x"D6",x"A9",x"80",x"85",x"2A",x"68",x"D0",x"D0", -- 0x1648
		x"A6",x"A6",x"A5",x"A7",x"86",x"A2",x"85",x"A3", -- 0x1650
		x"A0",x"00",x"84",x"BE",x"84",x"BD",x"A5",x"A0", -- 0x1658
		x"A6",x"A1",x"85",x"CE",x"86",x"CF",x"A9",x"88", -- 0x1660
		x"A2",x"00",x"85",x"91",x"86",x"92",x"C5",x"85", -- 0x1668
		x"F0",x"05",x"20",x"F1",x"D6",x"F0",x"F7",x"A9", -- 0x1670
		x"07",x"85",x"C2",x"A5",x"9C",x"A6",x"9D",x"85", -- 0x1678
		x"91",x"86",x"92",x"E4",x"9F",x"D0",x"04",x"C5", -- 0x1680
		x"9E",x"F0",x"05",x"20",x"E7",x"D6",x"F0",x"F3", -- 0x1688
		x"85",x"C7",x"86",x"C8",x"A9",x"03",x"85",x"C2", -- 0x1690
		x"A5",x"C7",x"A6",x"C8",x"E4",x"A1",x"D0",x"07", -- 0x1698
		x"C5",x"A0",x"D0",x"03",x"4C",x"30",x"D7",x"85", -- 0x16A0
		x"91",x"86",x"92",x"A0",x"00",x"B1",x"91",x"AA", -- 0x16A8
		x"C8",x"B1",x"91",x"08",x"C8",x"B1",x"91",x"65", -- 0x16B0
		x"C7",x"85",x"C7",x"C8",x"B1",x"91",x"65",x"C8", -- 0x16B8
		x"85",x"C8",x"28",x"10",x"D3",x"8A",x"30",x"D0", -- 0x16C0
		x"C8",x"B1",x"91",x"A0",x"00",x"0A",x"69",x"05", -- 0x16C8
		x"65",x"91",x"85",x"91",x"90",x"02",x"E6",x"92", -- 0x16D0
		x"A6",x"92",x"E4",x"C8",x"D0",x"04",x"C5",x"C7", -- 0x16D8
		x"F0",x"BA",x"20",x"F1",x"D6",x"F0",x"F3",x"B1", -- 0x16E0
		x"91",x"30",x"35",x"C8",x"B1",x"91",x"10",x"30", -- 0x16E8
		x"C8",x"B1",x"91",x"F0",x"2B",x"C8",x"B1",x"91", -- 0x16F0
		x"AA",x"C8",x"B1",x"91",x"C5",x"A3",x"90",x"06", -- 0x16F8
		x"D0",x"1E",x"E4",x"A2",x"B0",x"1A",x"C5",x"CF", -- 0x1700
		x"90",x"16",x"D0",x"04",x"E4",x"CE",x"90",x"10", -- 0x1708
		x"86",x"CE",x"85",x"CF",x"A5",x"91",x"A6",x"92", -- 0x1710
		x"85",x"BD",x"86",x"BE",x"A5",x"C2",x"85",x"C4", -- 0x1718
		x"A5",x"C2",x"18",x"65",x"91",x"85",x"91",x"90", -- 0x1720
		x"02",x"E6",x"92",x"A6",x"92",x"A0",x"00",x"60", -- 0x1728
		x"A5",x"BE",x"05",x"BD",x"F0",x"F5",x"A5",x"C4", -- 0x1730
		x"29",x"04",x"4A",x"A8",x"85",x"C4",x"B1",x"BD", -- 0x1738
		x"65",x"CE",x"85",x"C9",x"A5",x"CF",x"69",x"00", -- 0x1740
		x"85",x"CA",x"A5",x"A2",x"A6",x"A3",x"85",x"C7", -- 0x1748
		x"86",x"C8",x"20",x"FB",x"C3",x"A4",x"C4",x"C8", -- 0x1750
		x"A5",x"C7",x"91",x"BD",x"AA",x"E6",x"C8",x"A5", -- 0x1758
		x"C8",x"C8",x"91",x"BD",x"4C",x"54",x"D6",x"A5", -- 0x1760
		x"D4",x"48",x"A5",x"D3",x"48",x"20",x"00",x"D0", -- 0x1768
		x"20",x"08",x"CF",x"68",x"85",x"DE",x"68",x"85", -- 0x1770
		x"DF",x"A0",x"00",x"B1",x"DE",x"18",x"71",x"D3", -- 0x1778
		x"90",x"05",x"A2",x"B5",x"4C",x"7E",x"C4",x"20", -- 0x1780
		x"A3",x"D5",x"20",x"A4",x"D7",x"A5",x"BF",x"A4", -- 0x1788
		x"C0",x"20",x"D4",x"D7",x"20",x"B6",x"D7",x"A5", -- 0x1790
		x"DE",x"A4",x"DF",x"20",x"D4",x"D7",x"20",x"F4", -- 0x1798
		x"D5",x"4C",x"31",x"CF",x"A0",x"00",x"B1",x"DE", -- 0x17A0
		x"48",x"C8",x"B1",x"DE",x"AA",x"C8",x"B1",x"DE", -- 0x17A8
		x"A8",x"68",x"86",x"91",x"84",x"92",x"A8",x"F0", -- 0x17B0
		x"0A",x"48",x"88",x"B1",x"91",x"91",x"A4",x"98", -- 0x17B8
		x"D0",x"F8",x"68",x"18",x"65",x"A4",x"85",x"A4", -- 0x17C0
		x"90",x"02",x"E6",x"A5",x"60",x"20",x"08",x"CF", -- 0x17C8
		x"A5",x"D3",x"A4",x"D4",x"85",x"91",x"84",x"92", -- 0x17D0
		x"20",x"05",x"D8",x"08",x"A0",x"00",x"B1",x"91", -- 0x17D8
		x"48",x"C8",x"B1",x"91",x"AA",x"C8",x"B1",x"91", -- 0x17E0
		x"A8",x"68",x"28",x"D0",x"13",x"C4",x"A3",x"D0", -- 0x17E8
		x"0F",x"E4",x"A2",x"D0",x"0B",x"48",x"18",x"65", -- 0x17F0
		x"A2",x"85",x"A2",x"90",x"02",x"E6",x"A3",x"68", -- 0x17F8
		x"86",x"91",x"84",x"92",x"60",x"C4",x"87",x"D0", -- 0x1800
		x"0C",x"C5",x"86",x"D0",x"08",x"85",x"85",x"E9", -- 0x1808
		x"03",x"85",x"86",x"A0",x"00",x"60",x"20",x"CB", -- 0x1810
		x"D8",x"8A",x"48",x"A9",x"01",x"20",x"AB",x"D5", -- 0x1818
		x"68",x"A0",x"00",x"91",x"D1",x"68",x"68",x"4C", -- 0x1820
		x"F4",x"D5",x"20",x"8B",x"D8",x"D1",x"BF",x"98", -- 0x1828
		x"90",x"04",x"B1",x"BF",x"AA",x"98",x"48",x"8A", -- 0x1830
		x"48",x"20",x"AB",x"D5",x"A5",x"BF",x"A4",x"C0", -- 0x1838
		x"20",x"D4",x"D7",x"68",x"A8",x"68",x"18",x"65", -- 0x1840
		x"91",x"85",x"91",x"90",x"02",x"E6",x"92",x"98", -- 0x1848
		x"20",x"B6",x"D7",x"4C",x"F4",x"D5",x"20",x"8B", -- 0x1850
		x"D8",x"18",x"F1",x"BF",x"49",x"FF",x"4C",x"30", -- 0x1858
		x"D8",x"A9",x"FF",x"85",x"D4",x"20",x"E8",x"00", -- 0x1860
		x"C9",x"29",x"F0",x"06",x"20",x"65",x"D0",x"20", -- 0x1868
		x"C8",x"D8",x"20",x"8B",x"D8",x"F0",x"4B",x"CA", -- 0x1870
		x"8A",x"48",x"18",x"A2",x"00",x"F1",x"BF",x"B0", -- 0x1878
		x"B6",x"49",x"FF",x"C5",x"D4",x"90",x"B1",x"A5", -- 0x1880
		x"D4",x"B0",x"AD",x"20",x"5F",x"D0",x"68",x"A8", -- 0x1888
		x"68",x"85",x"C4",x"68",x"68",x"68",x"AA",x"68", -- 0x1890
		x"85",x"BF",x"68",x"85",x"C0",x"A5",x"C4",x"48", -- 0x1898
		x"98",x"48",x"A0",x"00",x"8A",x"60",x"20",x"AC", -- 0x18A0
		x"D8",x"4C",x"B6",x"D4",x"20",x"CD",x"D7",x"A2", -- 0x18A8
		x"00",x"86",x"28",x"A8",x"60",x"20",x"AC",x"D8", -- 0x18B0
		x"F0",x"08",x"A0",x"00",x"B1",x"91",x"A8",x"4C", -- 0x18B8
		x"B6",x"D4",x"4C",x"36",x"D3",x"20",x"E2",x"00", -- 0x18C0
		x"20",x"03",x"CF",x"20",x"A2",x"D2",x"A6",x"D3", -- 0x18C8
		x"D0",x"F0",x"A6",x"D4",x"4C",x"E8",x"00",x"20", -- 0x18D0
		x"AC",x"D8",x"D0",x"03",x"4C",x"B2",x"DB",x"A6", -- 0x18D8
		x"E9",x"A4",x"EA",x"86",x"E0",x"84",x"E1",x"A6", -- 0x18E0
		x"91",x"86",x"E9",x"18",x"65",x"91",x"85",x"93", -- 0x18E8
		x"A6",x"92",x"86",x"EA",x"90",x"01",x"E8",x"86", -- 0x18F0
		x"94",x"A0",x"00",x"B1",x"93",x"48",x"A9",x"00", -- 0x18F8
		x"91",x"93",x"20",x"E8",x"00",x"20",x"E7",x"DF", -- 0x1900
		x"68",x"A0",x"00",x"91",x"93",x"A6",x"E0",x"A4", -- 0x1908
		x"E1",x"86",x"E9",x"84",x"EA",x"60",x"20",x"03", -- 0x1910
		x"CF",x"20",x"22",x"D9",x"20",x"65",x"D0",x"4C", -- 0x1918
		x"C8",x"D8",x"A5",x"D5",x"30",x"9C",x"A5",x"D0", -- 0x1920
		x"C9",x"91",x"B0",x"96",x"20",x"8C",x"DF",x"A5", -- 0x1928
		x"D3",x"A4",x"D4",x"84",x"33",x"85",x"34",x"60", -- 0x1930
		x"A5",x"34",x"48",x"A5",x"33",x"48",x"20",x"22", -- 0x1938
		x"D9",x"A0",x"00",x"B1",x"33",x"A8",x"68",x"85", -- 0x1940
		x"33",x"68",x"85",x"34",x"4C",x"B6",x"D4",x"20", -- 0x1948
		x"16",x"D9",x"8A",x"A0",x"00",x"91",x"33",x"60", -- 0x1950
		x"20",x"03",x"CF",x"20",x"22",x"D9",x"A4",x"33", -- 0x1958
		x"A6",x"34",x"A9",x"02",x"4C",x"C9",x"EE",x"20", -- 0x1960
		x"53",x"E8",x"A5",x"33",x"A4",x"34",x"85",x"1D", -- 0x1968
		x"84",x"1E",x"20",x"65",x"D0",x"20",x"53",x"E8", -- 0x1970
		x"A0",x"01",x"B9",x"33",x"00",x"91",x"1D",x"88", -- 0x1978
		x"10",x"F8",x"60",x"20",x"22",x"D9",x"A0",x"01", -- 0x1980
		x"B1",x"33",x"48",x"88",x"B1",x"33",x"A8",x"68", -- 0x1988
		x"4C",x"40",x"DF",x"48",x"4A",x"4A",x"4A",x"4A", -- 0x1990
		x"20",x"9C",x"D9",x"68",x"29",x"0F",x"09",x"30", -- 0x1998
		x"C9",x"3A",x"90",x"02",x"69",x"06",x"C9",x"30", -- 0x19A0
		x"D0",x"04",x"A4",x"2F",x"F0",x"06",x"85",x"2F", -- 0x19A8
		x"9D",x"00",x"01",x"E8",x"60",x"20",x"22",x"D9", -- 0x19B0
		x"A2",x"00",x"86",x"2F",x"A9",x"23",x"85",x"FF", -- 0x19B8
		x"A5",x"34",x"20",x"93",x"D9",x"A5",x"33",x"20", -- 0x19C0
		x"93",x"D9",x"8A",x"D0",x"06",x"A9",x"30",x"9D", -- 0x19C8
		x"00",x"01",x"E8",x"A9",x"00",x"9D",x"00",x"01", -- 0x19D0
		x"4C",x"9B",x"D5",x"4C",x"70",x"D0",x"20",x"21", -- 0x19D8
		x"EC",x"20",x"C8",x"D8",x"8A",x"F0",x"06",x"CA", -- 0x19E0
		x"D0",x"F1",x"A9",x"09",x"2C",x"A9",x"08",x"A2", -- 0x19E8
		x"10",x"8E",x"F8",x"02",x"A2",x"1B",x"48",x"8A", -- 0x19F0
		x"20",x"0C",x"DA",x"AD",x"F8",x"02",x"A0",x"27", -- 0x19F8
		x"91",x"1F",x"88",x"D0",x"FB",x"68",x"91",x"1F", -- 0x1A00
		x"CA",x"D0",x"EB",x"60",x"20",x"31",x"F7",x"84", -- 0x1A08
		x"20",x"18",x"69",x"80",x"48",x"85",x"1F",x"A9", -- 0x1A10
		x"BB",x"65",x"20",x"85",x"20",x"68",x"60",x"4C", -- 0x1A18
		x"C2",x"D8",x"20",x"F6",x"DA",x"20",x"C8",x"D8", -- 0x1A20
		x"E0",x"28",x"B0",x"F3",x"8E",x"F8",x"02",x"20", -- 0x1A28
		x"65",x"D0",x"20",x"C8",x"D8",x"E0",x"1B",x"B0", -- 0x1A30
		x"E6",x"E8",x"8A",x"20",x"0C",x"DA",x"60",x"20", -- 0x1A38
		x"62",x"D0",x"20",x"22",x"DA",x"20",x"5F",x"D0", -- 0x1A40
		x"AC",x"F8",x"02",x"B1",x"1F",x"A8",x"4C",x"B6", -- 0x1A48
		x"D4",x"20",x"22",x"DA",x"20",x"65",x"D0",x"20", -- 0x1A50
		x"17",x"CF",x"24",x"28",x"10",x"1D",x"20",x"D0", -- 0x1A58
		x"D7",x"AA",x"18",x"AD",x"F8",x"02",x"65",x"1F", -- 0x1A60
		x"90",x"02",x"E6",x"20",x"85",x"1F",x"A0",x"00", -- 0x1A68
		x"E8",x"CA",x"F0",x"10",x"B1",x"91",x"91",x"1F", -- 0x1A70
		x"C8",x"D0",x"F6",x"20",x"CB",x"D8",x"8A",x"AC", -- 0x1A78
		x"F8",x"02",x"91",x"1F",x"60",x"D0",x"17",x"A9", -- 0x1A80
		x"03",x"20",x"37",x"C4",x"A5",x"EA",x"48",x"A5", -- 0x1A88
		x"E9",x"48",x"A5",x"A9",x"48",x"A5",x"A8",x"48", -- 0x1A90
		x"A9",x"8B",x"48",x"4C",x"C1",x"C8",x"4C",x"70", -- 0x1A98
		x"D0",x"A9",x"FF",x"85",x"B9",x"20",x"C6",x"C3", -- 0x1AA0
		x"9A",x"C9",x"8B",x"F0",x"05",x"A2",x"F5",x"4C", -- 0x1AA8
		x"7E",x"C4",x"C0",x"10",x"D0",x"05",x"84",x"D0", -- 0x1AB0
		x"98",x"D0",x"06",x"20",x"E8",x"00",x"20",x"17", -- 0x1AB8
		x"CF",x"68",x"A5",x"D0",x"F0",x"05",x"68",x"68", -- 0x1AC0
		x"68",x"68",x"60",x"68",x"85",x"A8",x"68",x"85", -- 0x1AC8
		x"A9",x"68",x"85",x"E9",x"68",x"85",x"EA",x"4C", -- 0x1AD0
		x"8C",x"DA",x"20",x"78",x"EB",x"08",x"48",x"10", -- 0x1AD8
		x"03",x"A9",x"01",x"2C",x"A9",x"00",x"20",x"AB", -- 0x1AE0
		x"D5",x"68",x"28",x"10",x"04",x"A0",x"00",x"91", -- 0x1AE8
		x"D1",x"68",x"68",x"4C",x"F4",x"D5",x"AD",x"C0", -- 0x1AF0
		x"02",x"29",x"01",x"F0",x"05",x"A2",x"A3",x"4C", -- 0x1AF8
		x"7E",x"C4",x"60",x"60",x"A9",x"05",x"A0",x"E2", -- 0x1B00
		x"4C",x"22",x"DB",x"20",x"51",x"DD",x"A5",x"D5", -- 0x1B08
		x"49",x"FF",x"85",x"D5",x"45",x"DD",x"85",x"DE", -- 0x1B10
		x"A5",x"D0",x"4C",x"25",x"DB",x"20",x"54",x"DC", -- 0x1B18
		x"90",x"3C",x"20",x"51",x"DD",x"D0",x"03",x"4C", -- 0x1B20
		x"D5",x"DE",x"A6",x"DF",x"86",x"C5",x"A2",x"D8", -- 0x1B28
		x"A5",x"D8",x"A8",x"F0",x"CE",x"38",x"E5",x"D0", -- 0x1B30
		x"F0",x"24",x"90",x"12",x"84",x"D0",x"A4",x"DD", -- 0x1B38
		x"84",x"D5",x"49",x"FF",x"69",x"00",x"A0",x"00", -- 0x1B40
		x"84",x"C5",x"A2",x"D0",x"D0",x"04",x"A0",x"00", -- 0x1B48
		x"84",x"DF",x"C9",x"F9",x"30",x"C7",x"A8",x"A5", -- 0x1B50
		x"DF",x"56",x"01",x"20",x"6B",x"DC",x"24",x"DE", -- 0x1B58
		x"10",x"57",x"A0",x"D0",x"E0",x"D8",x"F0",x"02", -- 0x1B60
		x"A0",x"D8",x"38",x"49",x"FF",x"65",x"C5",x"85", -- 0x1B68
		x"DF",x"B9",x"04",x"00",x"F5",x"04",x"85",x"D4", -- 0x1B70
		x"B9",x"03",x"00",x"F5",x"03",x"85",x"D3",x"B9", -- 0x1B78
		x"02",x"00",x"F5",x"02",x"85",x"D2",x"B9",x"01", -- 0x1B80
		x"00",x"F5",x"01",x"85",x"D1",x"B0",x"03",x"20", -- 0x1B88
		x"02",x"DC",x"A0",x"00",x"98",x"18",x"A6",x"D1", -- 0x1B90
		x"D0",x"4A",x"A6",x"D2",x"86",x"D1",x"A6",x"D3", -- 0x1B98
		x"86",x"D2",x"A6",x"D4",x"86",x"D3",x"A6",x"DF", -- 0x1BA0
		x"86",x"D4",x"84",x"DF",x"69",x"08",x"C9",x"28", -- 0x1BA8
		x"D0",x"E4",x"A9",x"00",x"85",x"D0",x"85",x"D5", -- 0x1BB0
		x"60",x"65",x"C5",x"85",x"DF",x"A5",x"D4",x"65", -- 0x1BB8
		x"DC",x"85",x"D4",x"A5",x"D3",x"65",x"DB",x"85", -- 0x1BC0
		x"D3",x"A5",x"D2",x"65",x"DA",x"85",x"D2",x"A5", -- 0x1BC8
		x"D1",x"65",x"D9",x"85",x"D1",x"4C",x"F1",x"DB", -- 0x1BD0
		x"69",x"01",x"06",x"DF",x"26",x"D4",x"26",x"D3", -- 0x1BD8
		x"26",x"D2",x"26",x"D1",x"10",x"F2",x"38",x"E5", -- 0x1BE0
		x"D0",x"B0",x"C7",x"49",x"FF",x"69",x"01",x"85", -- 0x1BE8
		x"D0",x"90",x"0E",x"E6",x"D0",x"F0",x"42",x"66", -- 0x1BF0
		x"D1",x"66",x"D2",x"66",x"D3",x"66",x"D4",x"66", -- 0x1BF8
		x"DF",x"60",x"A5",x"D5",x"49",x"FF",x"85",x"D5", -- 0x1C00
		x"A5",x"D1",x"49",x"FF",x"85",x"D1",x"A5",x"D2", -- 0x1C08
		x"49",x"FF",x"85",x"D2",x"A5",x"D3",x"49",x"FF", -- 0x1C10
		x"85",x"D3",x"A5",x"D4",x"49",x"FF",x"85",x"D4", -- 0x1C18
		x"A5",x"DF",x"49",x"FF",x"85",x"DF",x"E6",x"DF", -- 0x1C20
		x"D0",x"0E",x"E6",x"D4",x"D0",x"0A",x"E6",x"D3", -- 0x1C28
		x"D0",x"06",x"E6",x"D2",x"D0",x"02",x"E6",x"D1", -- 0x1C30
		x"60",x"A2",x"45",x"4C",x"7E",x"C4",x"A2",x"94", -- 0x1C38
		x"B4",x"04",x"84",x"DF",x"B4",x"03",x"94",x"04", -- 0x1C40
		x"B4",x"02",x"94",x"03",x"B4",x"01",x"94",x"02", -- 0x1C48
		x"A4",x"D7",x"94",x"01",x"69",x"08",x"30",x"E8", -- 0x1C50
		x"F0",x"E6",x"E9",x"08",x"A8",x"A5",x"DF",x"B0", -- 0x1C58
		x"14",x"16",x"01",x"90",x"02",x"F6",x"01",x"76", -- 0x1C60
		x"01",x"76",x"01",x"76",x"02",x"76",x"03",x"76", -- 0x1C68
		x"04",x"6A",x"C8",x"D0",x"EC",x"18",x"60",x"82", -- 0x1C70
		x"13",x"5D",x"8D",x"DE",x"82",x"49",x"0F",x"DA", -- 0x1C78
		x"9E",x"81",x"00",x"00",x"00",x"00",x"03",x"7F", -- 0x1C80
		x"5E",x"56",x"CB",x"79",x"80",x"13",x"9B",x"0B", -- 0x1C88
		x"64",x"80",x"76",x"38",x"93",x"16",x"82",x"38", -- 0x1C90
		x"AA",x"3B",x"20",x"80",x"35",x"04",x"F3",x"34", -- 0x1C98
		x"81",x"35",x"04",x"F3",x"34",x"80",x"80",x"00", -- 0x1CA0
		x"00",x"00",x"80",x"31",x"72",x"17",x"F8",x"20", -- 0x1CA8
		x"13",x"DF",x"F0",x"02",x"10",x"03",x"4C",x"36", -- 0x1CB0
		x"D3",x"A5",x"D0",x"E9",x"7F",x"48",x"A9",x"80", -- 0x1CB8
		x"85",x"D0",x"A9",x"9B",x"A0",x"DC",x"20",x"22", -- 0x1CC0
		x"DB",x"A9",x"A0",x"A0",x"DC",x"20",x"E4",x"DD", -- 0x1CC8
		x"A9",x"81",x"A0",x"DC",x"20",x"0B",x"DB",x"A9", -- 0x1CD0
		x"86",x"A0",x"DC",x"20",x"FD",x"E2",x"A9",x"A5", -- 0x1CD8
		x"A0",x"DC",x"20",x"22",x"DB",x"68",x"20",x"76", -- 0x1CE0
		x"E0",x"A9",x"AA",x"A0",x"DC",x"20",x"51",x"DD", -- 0x1CE8
		x"D0",x"03",x"4C",x"50",x"DD",x"20",x"7C",x"DD", -- 0x1CF0
		x"A9",x"00",x"85",x"95",x"85",x"96",x"85",x"97", -- 0x1CF8
		x"85",x"98",x"A5",x"DF",x"20",x"1E",x"DD",x"A5", -- 0x1D00
		x"D4",x"20",x"1E",x"DD",x"A5",x"D3",x"20",x"1E", -- 0x1D08
		x"DD",x"A5",x"D2",x"20",x"1E",x"DD",x"A5",x"D1", -- 0x1D10
		x"20",x"23",x"DD",x"4C",x"64",x"DE",x"D0",x"03", -- 0x1D18
		x"4C",x"3E",x"DC",x"4A",x"09",x"80",x"A8",x"90", -- 0x1D20
		x"19",x"18",x"A5",x"98",x"65",x"DC",x"85",x"98", -- 0x1D28
		x"A5",x"97",x"65",x"DB",x"85",x"97",x"A5",x"96", -- 0x1D30
		x"65",x"DA",x"85",x"96",x"A5",x"95",x"65",x"D9", -- 0x1D38
		x"85",x"95",x"66",x"95",x"66",x"96",x"66",x"97", -- 0x1D40
		x"66",x"98",x"66",x"DF",x"98",x"4A",x"D0",x"D6", -- 0x1D48
		x"60",x"85",x"91",x"84",x"92",x"A0",x"04",x"B1", -- 0x1D50
		x"91",x"85",x"DC",x"88",x"B1",x"91",x"85",x"DB", -- 0x1D58
		x"88",x"B1",x"91",x"85",x"DA",x"88",x"B1",x"91", -- 0x1D60
		x"85",x"DD",x"45",x"D5",x"85",x"DE",x"A5",x"DD", -- 0x1D68
		x"09",x"80",x"85",x"D9",x"88",x"B1",x"91",x"85", -- 0x1D70
		x"D8",x"A5",x"D0",x"60",x"A5",x"D8",x"F0",x"1F", -- 0x1D78
		x"18",x"65",x"D0",x"90",x"04",x"30",x"1D",x"18", -- 0x1D80
		x"2C",x"10",x"14",x"69",x"80",x"85",x"D0",x"D0", -- 0x1D88
		x"03",x"4C",x"B6",x"DB",x"A5",x"DE",x"85",x"D5", -- 0x1D90
		x"60",x"A5",x"D5",x"49",x"FF",x"30",x"05",x"68", -- 0x1D98
		x"68",x"4C",x"B2",x"DB",x"4C",x"39",x"DC",x"20", -- 0x1DA0
		x"E5",x"DE",x"AA",x"F0",x"10",x"18",x"69",x"02", -- 0x1DA8
		x"B0",x"F2",x"A2",x"00",x"86",x"DE",x"20",x"32", -- 0x1DB0
		x"DB",x"E6",x"D0",x"F0",x"E7",x"60",x"84",x"20", -- 0x1DB8
		x"00",x"00",x"00",x"20",x"E5",x"DE",x"A9",x"BE", -- 0x1DC0
		x"A0",x"DD",x"A2",x"00",x"86",x"DE",x"20",x"7B", -- 0x1DC8
		x"DE",x"4C",x"E7",x"DD",x"20",x"AF",x"DC",x"20", -- 0x1DD0
		x"E5",x"DE",x"A9",x"77",x"A0",x"DC",x"20",x"7B", -- 0x1DD8
		x"DE",x"4C",x"E7",x"DD",x"20",x"51",x"DD",x"F0", -- 0x1DE0
		x"76",x"20",x"F4",x"DE",x"A9",x"00",x"38",x"E5", -- 0x1DE8
		x"D0",x"85",x"D0",x"20",x"7C",x"DD",x"E6",x"D0", -- 0x1DF0
		x"F0",x"AA",x"A2",x"FC",x"A9",x"01",x"A4",x"D9", -- 0x1DF8
		x"C4",x"D1",x"D0",x"10",x"A4",x"DA",x"C4",x"D2", -- 0x1E00
		x"D0",x"0A",x"A4",x"DB",x"C4",x"D3",x"D0",x"04", -- 0x1E08
		x"A4",x"DC",x"C4",x"D4",x"08",x"2A",x"90",x"09", -- 0x1E10
		x"E8",x"95",x"98",x"F0",x"32",x"10",x"34",x"A9", -- 0x1E18
		x"01",x"28",x"B0",x"0E",x"06",x"DC",x"26",x"DB", -- 0x1E20
		x"26",x"DA",x"26",x"D9",x"B0",x"E6",x"30",x"CE", -- 0x1E28
		x"10",x"E2",x"A8",x"A5",x"DC",x"E5",x"D4",x"85", -- 0x1E30
		x"DC",x"A5",x"DB",x"E5",x"D3",x"85",x"DB",x"A5", -- 0x1E38
		x"DA",x"E5",x"D2",x"85",x"DA",x"A5",x"D9",x"E5", -- 0x1E40
		x"D1",x"85",x"D9",x"98",x"4C",x"24",x"DE",x"A9", -- 0x1E48
		x"40",x"D0",x"CE",x"0A",x"0A",x"0A",x"0A",x"0A", -- 0x1E50
		x"0A",x"85",x"DF",x"28",x"4C",x"64",x"DE",x"A2", -- 0x1E58
		x"85",x"4C",x"7E",x"C4",x"A5",x"95",x"85",x"D1", -- 0x1E60
		x"A5",x"96",x"85",x"D2",x"A5",x"97",x"85",x"D3", -- 0x1E68
		x"A5",x"98",x"85",x"D4",x"4C",x"92",x"DB",x"A9", -- 0x1E70
		x"7C",x"A0",x"DC",x"85",x"91",x"84",x"92",x"A0", -- 0x1E78
		x"04",x"B1",x"91",x"85",x"D4",x"88",x"B1",x"91", -- 0x1E80
		x"85",x"D3",x"88",x"B1",x"91",x"85",x"D2",x"88", -- 0x1E88
		x"B1",x"91",x"85",x"D5",x"09",x"80",x"85",x"D1", -- 0x1E90
		x"88",x"B1",x"91",x"85",x"D0",x"84",x"DF",x"60", -- 0x1E98
		x"A2",x"CB",x"2C",x"A2",x"C6",x"A0",x"00",x"F0", -- 0x1EA0
		x"04",x"A6",x"B8",x"A4",x"B9",x"20",x"F4",x"DE", -- 0x1EA8
		x"86",x"91",x"84",x"92",x"A0",x"04",x"A5",x"D4", -- 0x1EB0
		x"91",x"91",x"88",x"A5",x"D3",x"91",x"91",x"88", -- 0x1EB8
		x"A5",x"D2",x"91",x"91",x"88",x"A5",x"D5",x"09", -- 0x1EC0
		x"7F",x"25",x"D1",x"91",x"91",x"88",x"A5",x"D0", -- 0x1EC8
		x"91",x"91",x"84",x"DF",x"60",x"A5",x"DD",x"85", -- 0x1ED0
		x"D5",x"A2",x"05",x"B5",x"D7",x"95",x"CF",x"CA", -- 0x1ED8
		x"D0",x"F9",x"86",x"DF",x"60",x"20",x"F4",x"DE", -- 0x1EE0
		x"A2",x"06",x"B5",x"CF",x"95",x"D7",x"CA",x"D0", -- 0x1EE8
		x"F9",x"86",x"DF",x"60",x"A5",x"D0",x"F0",x"FB", -- 0x1EF0
		x"06",x"DF",x"90",x"F7",x"20",x"2A",x"DC",x"D0", -- 0x1EF8
		x"F2",x"4C",x"F3",x"DB",x"20",x"A9",x"D2",x"46", -- 0x1F00
		x"D4",x"B0",x"04",x"A9",x"00",x"F0",x"15",x"A9", -- 0x1F08
		x"FF",x"30",x"11",x"A5",x"D0",x"F0",x"09",x"A5", -- 0x1F10
		x"D5",x"2A",x"A9",x"FF",x"B0",x"02",x"A9",x"01", -- 0x1F18
		x"60",x"20",x"13",x"DF",x"85",x"D1",x"A9",x"00", -- 0x1F20
		x"85",x"D2",x"A2",x"88",x"A5",x"D1",x"49",x"FF", -- 0x1F28
		x"2A",x"A9",x"00",x"85",x"D4",x"85",x"D3",x"86", -- 0x1F30
		x"D0",x"85",x"DF",x"85",x"D5",x"4C",x"8D",x"DB", -- 0x1F38
		x"85",x"D1",x"84",x"D2",x"A2",x"90",x"38",x"B0", -- 0x1F40
		x"E8",x"46",x"D5",x"60",x"85",x"93",x"84",x"94", -- 0x1F48
		x"A0",x"00",x"B1",x"93",x"C8",x"AA",x"F0",x"BB", -- 0x1F50
		x"B1",x"93",x"45",x"D5",x"30",x"B9",x"E4",x"D0", -- 0x1F58
		x"D0",x"21",x"B1",x"93",x"09",x"80",x"C5",x"D1", -- 0x1F60
		x"D0",x"19",x"C8",x"B1",x"93",x"C5",x"D2",x"D0", -- 0x1F68
		x"12",x"C8",x"B1",x"93",x"C5",x"D3",x"D0",x"0B", -- 0x1F70
		x"C8",x"A9",x"7F",x"C5",x"DF",x"B1",x"93",x"E5", -- 0x1F78
		x"D4",x"F0",x"28",x"A5",x"D5",x"90",x"02",x"49", -- 0x1F80
		x"FF",x"4C",x"19",x"DF",x"A5",x"D0",x"F0",x"4A", -- 0x1F88
		x"38",x"E9",x"A0",x"24",x"D5",x"10",x"09",x"AA", -- 0x1F90
		x"A9",x"FF",x"85",x"D7",x"20",x"08",x"DC",x"8A", -- 0x1F98
		x"A2",x"D0",x"C9",x"F9",x"10",x"06",x"20",x"54", -- 0x1FA0
		x"DC",x"84",x"D7",x"60",x"A8",x"A5",x"D5",x"29", -- 0x1FA8
		x"80",x"46",x"D1",x"05",x"D1",x"85",x"D1",x"20", -- 0x1FB0
		x"6B",x"DC",x"84",x"D7",x"60",x"A5",x"D0",x"C9", -- 0x1FB8
		x"A0",x"B0",x"20",x"20",x"8C",x"DF",x"84",x"DF", -- 0x1FC0
		x"A5",x"D5",x"84",x"D5",x"49",x"80",x"2A",x"A9", -- 0x1FC8
		x"A0",x"85",x"D0",x"A5",x"D4",x"85",x"24",x"4C", -- 0x1FD0
		x"8D",x"DB",x"85",x"D1",x"85",x"D2",x"85",x"D3", -- 0x1FD8
		x"85",x"D4",x"A8",x"60",x"4C",x"81",x"E9",x"A0", -- 0x1FE0
		x"00",x"A2",x"0A",x"94",x"CC",x"CA",x"10",x"FB", -- 0x1FE8
		x"90",x"13",x"C9",x"23",x"F0",x"EE",x"C9",x"2D", -- 0x1FF0
		x"D0",x"04",x"86",x"D6",x"F0",x"04",x"C9",x"2B", -- 0x1FF8
		x"D0",x"05",x"20",x"E2",x"00",x"90",x"5B",x"C9", -- 0x2000
		x"2E",x"F0",x"2E",x"C9",x"45",x"D0",x"30",x"20", -- 0x2008
		x"E2",x"00",x"90",x"17",x"C9",x"CD",x"F0",x"0E", -- 0x2010
		x"C9",x"2D",x"F0",x"0A",x"C9",x"CC",x"F0",x"08", -- 0x2018
		x"C9",x"2B",x"F0",x"04",x"D0",x"07",x"66",x"CF", -- 0x2020
		x"20",x"E2",x"00",x"90",x"5C",x"24",x"CF",x"10", -- 0x2028
		x"0E",x"A9",x"00",x"38",x"E5",x"CD",x"4C",x"41", -- 0x2030
		x"E0",x"66",x"CE",x"24",x"CE",x"50",x"C3",x"A5", -- 0x2038
		x"CD",x"38",x"E5",x"CC",x"85",x"CD",x"F0",x"12", -- 0x2040
		x"10",x"09",x"20",x"C3",x"DD",x"E6",x"CD",x"D0", -- 0x2048
		x"F9",x"F0",x"07",x"20",x"A7",x"DD",x"C6",x"CD", -- 0x2050
		x"D0",x"F9",x"A5",x"D6",x"30",x"01",x"60",x"4C", -- 0x2058
		x"71",x"E2",x"48",x"24",x"CE",x"10",x"02",x"E6", -- 0x2060
		x"CC",x"20",x"A7",x"DD",x"68",x"38",x"E9",x"30", -- 0x2068
		x"20",x"76",x"E0",x"4C",x"02",x"E0",x"48",x"20", -- 0x2070
		x"E5",x"DE",x"68",x"20",x"24",x"DF",x"A5",x"DD", -- 0x2078
		x"45",x"D5",x"85",x"DE",x"A6",x"D0",x"4C",x"25", -- 0x2080
		x"DB",x"A5",x"CD",x"C9",x"0A",x"90",x"09",x"A9", -- 0x2088
		x"64",x"24",x"CF",x"30",x"11",x"4C",x"39",x"DC", -- 0x2090
		x"0A",x"0A",x"18",x"65",x"CD",x"0A",x"18",x"A0", -- 0x2098
		x"00",x"71",x"E9",x"38",x"E9",x"30",x"85",x"CD", -- 0x20A0
		x"4C",x"28",x"E0",x"9B",x"3E",x"BC",x"1F",x"FD", -- 0x20A8
		x"9E",x"6E",x"6B",x"27",x"FD",x"9E",x"6E",x"6B", -- 0x20B0
		x"28",x"00",x"A9",x"AD",x"A0",x"C3",x"20",x"D2", -- 0x20B8
		x"E0",x"A5",x"A9",x"A6",x"A8",x"85",x"D1",x"86", -- 0x20C0
		x"D2",x"A2",x"90",x"38",x"20",x"31",x"DF",x"20", -- 0x20C8
		x"D5",x"E0",x"4C",x"B0",x"CC",x"A0",x"01",x"A9", -- 0x20D0
		x"20",x"24",x"D5",x"10",x"02",x"A9",x"2D",x"99", -- 0x20D8
		x"FF",x"00",x"85",x"D5",x"84",x"E0",x"C8",x"A9", -- 0x20E0
		x"30",x"A6",x"D0",x"D0",x"03",x"4C",x"F8",x"E1", -- 0x20E8
		x"A9",x"00",x"E0",x"80",x"F0",x"02",x"B0",x"09", -- 0x20F0
		x"A9",x"B5",x"A0",x"E0",x"20",x"ED",x"DC",x"A9", -- 0x20F8
		x"F7",x"85",x"CC",x"A9",x"B0",x"A0",x"E0",x"20", -- 0x2100
		x"4C",x"DF",x"F0",x"1E",x"10",x"12",x"A9",x"AB", -- 0x2108
		x"A0",x"E0",x"20",x"4C",x"DF",x"F0",x"02",x"10", -- 0x2110
		x"0E",x"20",x"A7",x"DD",x"C6",x"CC",x"D0",x"EE", -- 0x2118
		x"20",x"C3",x"DD",x"E6",x"CC",x"D0",x"DC",x"20", -- 0x2120
		x"04",x"DB",x"20",x"8C",x"DF",x"A2",x"01",x"A5", -- 0x2128
		x"CC",x"18",x"69",x"0A",x"30",x"09",x"C9",x"0B", -- 0x2130
		x"B0",x"06",x"69",x"FF",x"AA",x"A9",x"02",x"38", -- 0x2138
		x"E9",x"02",x"85",x"CD",x"86",x"CC",x"8A",x"F0", -- 0x2140
		x"02",x"10",x"13",x"A4",x"E0",x"A9",x"2E",x"C8", -- 0x2148
		x"99",x"FF",x"00",x"8A",x"F0",x"06",x"A9",x"30", -- 0x2150
		x"C8",x"99",x"FF",x"00",x"84",x"E0",x"A0",x"00", -- 0x2158
		x"A2",x"80",x"A5",x"D4",x"18",x"79",x"0D",x"E2", -- 0x2160
		x"85",x"D4",x"A5",x"D3",x"79",x"0C",x"E2",x"85", -- 0x2168
		x"D3",x"A5",x"D2",x"79",x"0B",x"E2",x"85",x"D2", -- 0x2170
		x"A5",x"D1",x"79",x"0A",x"E2",x"85",x"D1",x"E8", -- 0x2178
		x"B0",x"04",x"10",x"DE",x"30",x"02",x"30",x"DA", -- 0x2180
		x"8A",x"90",x"04",x"49",x"FF",x"69",x"0A",x"69", -- 0x2188
		x"2F",x"C8",x"C8",x"C8",x"C8",x"84",x"B6",x"A4", -- 0x2190
		x"E0",x"C8",x"AA",x"29",x"7F",x"99",x"FF",x"00", -- 0x2198
		x"C6",x"CC",x"D0",x"06",x"A9",x"2E",x"C8",x"99", -- 0x21A0
		x"FF",x"00",x"84",x"E0",x"A4",x"B6",x"8A",x"49", -- 0x21A8
		x"FF",x"29",x"80",x"AA",x"C0",x"24",x"D0",x"AA", -- 0x21B0
		x"A4",x"E0",x"B9",x"FF",x"00",x"88",x"C9",x"30", -- 0x21B8
		x"F0",x"F8",x"C9",x"2E",x"F0",x"01",x"C8",x"A9", -- 0x21C0
		x"2B",x"A6",x"CD",x"F0",x"2E",x"10",x"08",x"A9", -- 0x21C8
		x"00",x"38",x"E5",x"CD",x"AA",x"A9",x"2D",x"99", -- 0x21D0
		x"01",x"01",x"A9",x"45",x"99",x"00",x"01",x"8A", -- 0x21D8
		x"A2",x"2F",x"38",x"E8",x"E9",x"0A",x"B0",x"FB", -- 0x21E0
		x"69",x"3A",x"99",x"03",x"01",x"8A",x"99",x"02", -- 0x21E8
		x"01",x"A9",x"00",x"99",x"04",x"01",x"F0",x"08", -- 0x21F0
		x"99",x"FF",x"00",x"A9",x"00",x"99",x"00",x"01", -- 0x21F8
		x"A9",x"00",x"A0",x"01",x"60",x"80",x"00",x"00", -- 0x2200
		x"00",x"00",x"FA",x"0A",x"1F",x"00",x"00",x"98", -- 0x2208
		x"96",x"80",x"FF",x"F0",x"BD",x"C0",x"00",x"01", -- 0x2210
		x"86",x"A0",x"FF",x"FF",x"D8",x"F0",x"00",x"00", -- 0x2218
		x"03",x"E8",x"FF",x"FF",x"FF",x"9C",x"00",x"00", -- 0x2220
		x"00",x"0A",x"FF",x"FF",x"FF",x"FF",x"20",x"E5", -- 0x2228
		x"DE",x"A9",x"05",x"A0",x"E2",x"20",x"7B",x"DE", -- 0x2230
		x"F0",x"70",x"A5",x"D8",x"D0",x"03",x"4C",x"B4", -- 0x2238
		x"DB",x"A2",x"BD",x"A0",x"00",x"20",x"AD",x"DE", -- 0x2240
		x"A5",x"DD",x"10",x"0F",x"20",x"BD",x"DF",x"A9", -- 0x2248
		x"BD",x"A0",x"00",x"20",x"4C",x"DF",x"D0",x"03", -- 0x2250
		x"98",x"A4",x"24",x"20",x"D7",x"DE",x"98",x"48", -- 0x2258
		x"20",x"AF",x"DC",x"A9",x"BD",x"A0",x"00",x"20", -- 0x2260
		x"ED",x"DC",x"20",x"AA",x"E2",x"68",x"4A",x"90", -- 0x2268
		x"0A",x"A5",x"D0",x"F0",x"06",x"A5",x"D5",x"49", -- 0x2270
		x"FF",x"85",x"D5",x"60",x"81",x"38",x"AA",x"3B", -- 0x2278
		x"29",x"07",x"71",x"34",x"58",x"3E",x"56",x"74", -- 0x2280
		x"16",x"7E",x"B3",x"1B",x"77",x"2F",x"EE",x"E3", -- 0x2288
		x"85",x"7A",x"1D",x"84",x"1C",x"2A",x"7C",x"63", -- 0x2290
		x"59",x"58",x"0A",x"7E",x"75",x"FD",x"E7",x"C6", -- 0x2298
		x"80",x"31",x"72",x"18",x"10",x"81",x"00",x"00", -- 0x22A0
		x"00",x"00",x"A9",x"7C",x"A0",x"E2",x"20",x"ED", -- 0x22A8
		x"DC",x"A5",x"DF",x"69",x"50",x"90",x"03",x"20", -- 0x22B0
		x"FC",x"DE",x"85",x"C5",x"20",x"E8",x"DE",x"A5", -- 0x22B8
		x"D0",x"C9",x"88",x"90",x"03",x"20",x"99",x"DD", -- 0x22C0
		x"20",x"BD",x"DF",x"A5",x"24",x"18",x"69",x"81", -- 0x22C8
		x"F0",x"F3",x"38",x"E9",x"01",x"48",x"A2",x"05", -- 0x22D0
		x"B5",x"D8",x"B4",x"D0",x"95",x"D0",x"94",x"D8", -- 0x22D8
		x"CA",x"10",x"F5",x"A5",x"C5",x"85",x"DF",x"20", -- 0x22E0
		x"0E",x"DB",x"20",x"71",x"E2",x"A9",x"81",x"A0", -- 0x22E8
		x"E2",x"20",x"13",x"E3",x"A9",x"00",x"85",x"DE", -- 0x22F0
		x"68",x"20",x"7E",x"DD",x"60",x"85",x"E0",x"84", -- 0x22F8
		x"E1",x"20",x"A3",x"DE",x"A9",x"C6",x"20",x"ED", -- 0x2300
		x"DC",x"20",x"17",x"E3",x"A9",x"C6",x"A0",x"00", -- 0x2308
		x"4C",x"ED",x"DC",x"85",x"E0",x"84",x"E1",x"20", -- 0x2310
		x"A0",x"DE",x"B1",x"E0",x"85",x"D6",x"A4",x"E0", -- 0x2318
		x"C8",x"98",x"D0",x"02",x"E6",x"E1",x"85",x"E0", -- 0x2320
		x"A4",x"E1",x"20",x"ED",x"DC",x"A5",x"E0",x"A4", -- 0x2328
		x"E1",x"18",x"69",x"05",x"90",x"01",x"C8",x"85", -- 0x2330
		x"E0",x"84",x"E1",x"20",x"22",x"DB",x"A9",x"CB", -- 0x2338
		x"A0",x"00",x"C6",x"D6",x"D0",x"E4",x"60",x"98", -- 0x2340
		x"35",x"44",x"7A",x"68",x"28",x"B1",x"46",x"20", -- 0x2348
		x"13",x"DF",x"AA",x"30",x"18",x"A9",x"FA",x"A0", -- 0x2350
		x"00",x"20",x"7B",x"DE",x"8A",x"F0",x"E7",x"A9", -- 0x2358
		x"47",x"A0",x"E3",x"20",x"ED",x"DC",x"A9",x"4B", -- 0x2360
		x"A0",x"E3",x"20",x"22",x"DB",x"A6",x"D4",x"A5", -- 0x2368
		x"D1",x"85",x"D4",x"86",x"D1",x"A9",x"00",x"85", -- 0x2370
		x"D5",x"A5",x"D0",x"85",x"DF",x"A9",x"80",x"85", -- 0x2378
		x"D0",x"20",x"92",x"DB",x"A2",x"FA",x"A0",x"00", -- 0x2380
		x"4C",x"AD",x"DE",x"A9",x"07",x"A0",x"E4",x"20", -- 0x2388
		x"22",x"DB",x"20",x"E5",x"DE",x"A9",x"0C",x"A0", -- 0x2390
		x"E4",x"A6",x"DD",x"20",x"CC",x"DD",x"20",x"E5", -- 0x2398
		x"DE",x"20",x"BD",x"DF",x"A9",x"00",x"85",x"DE", -- 0x23A0
		x"20",x"0E",x"DB",x"A9",x"11",x"A0",x"E4",x"20", -- 0x23A8
		x"0B",x"DB",x"A5",x"D5",x"48",x"10",x"0D",x"20", -- 0x23B0
		x"04",x"DB",x"A5",x"D5",x"30",x"09",x"A5",x"2D", -- 0x23B8
		x"49",x"FF",x"85",x"2D",x"20",x"71",x"E2",x"A9", -- 0x23C0
		x"11",x"A0",x"E4",x"20",x"22",x"DB",x"68",x"10", -- 0x23C8
		x"03",x"20",x"71",x"E2",x"A9",x"16",x"A0",x"E4", -- 0x23D0
		x"4C",x"FD",x"E2",x"20",x"A3",x"DE",x"A9",x"00", -- 0x23D8
		x"85",x"2D",x"20",x"92",x"E3",x"A2",x"BD",x"A0", -- 0x23E0
		x"00",x"20",x"88",x"E3",x"A9",x"C6",x"A0",x"00", -- 0x23E8
		x"20",x"7B",x"DE",x"A9",x"00",x"85",x"D5",x"A5", -- 0x23F0
		x"2D",x"20",x"03",x"E4",x"A9",x"BD",x"A0",x"00", -- 0x23F8
		x"4C",x"E4",x"DD",x"48",x"4C",x"C4",x"E3",x"81", -- 0x2400
		x"49",x"0F",x"DA",x"A2",x"83",x"49",x"0F",x"DA", -- 0x2408
		x"A2",x"7F",x"00",x"00",x"00",x"00",x"05",x"84", -- 0x2410
		x"E6",x"1A",x"2D",x"1B",x"86",x"28",x"07",x"FB", -- 0x2418
		x"F8",x"87",x"99",x"68",x"89",x"01",x"87",x"23", -- 0x2420
		x"35",x"DF",x"E1",x"86",x"A5",x"5D",x"E7",x"28", -- 0x2428
		x"83",x"49",x"0F",x"DA",x"A2",x"A1",x"54",x"46", -- 0x2430
		x"8F",x"13",x"8F",x"52",x"43",x"89",x"CD",x"A5", -- 0x2438
		x"D5",x"48",x"10",x"03",x"20",x"71",x"E2",x"A5", -- 0x2440
		x"D0",x"48",x"C9",x"81",x"90",x"07",x"A9",x"81", -- 0x2448
		x"A0",x"DC",x"20",x"E4",x"DD",x"A9",x"6F",x"A0", -- 0x2450
		x"E4",x"20",x"FD",x"E2",x"68",x"C9",x"81",x"90", -- 0x2458
		x"07",x"A9",x"07",x"A0",x"E4",x"20",x"0B",x"DB", -- 0x2460
		x"68",x"10",x"03",x"4C",x"71",x"E2",x"60",x"0B", -- 0x2468
		x"76",x"B3",x"83",x"BD",x"D3",x"79",x"1E",x"F4", -- 0x2470
		x"A6",x"F5",x"7B",x"83",x"FC",x"B0",x"10",x"7C", -- 0x2478
		x"0C",x"1F",x"67",x"CA",x"7C",x"DE",x"53",x"CB", -- 0x2480
		x"C1",x"7D",x"14",x"64",x"70",x"4C",x"7D",x"B7", -- 0x2488
		x"EA",x"51",x"7A",x"7D",x"63",x"30",x"88",x"7E", -- 0x2490
		x"7E",x"92",x"44",x"99",x"3A",x"7E",x"4C",x"CC", -- 0x2498
		x"91",x"C7",x"7F",x"AA",x"AA",x"AA",x"13",x"81", -- 0x24A0
		x"00",x"00",x"00",x"00",x"20",x"35",x"E7",x"20", -- 0x24A8
		x"C9",x"E6",x"C9",x"24",x"D0",x"F9",x"8E",x"B1", -- 0x24B0
		x"02",x"A2",x"09",x"20",x"C9",x"E6",x"9D",x"A7", -- 0x24B8
		x"02",x"CA",x"D0",x"F7",x"20",x"C9",x"E6",x"F0", -- 0x24C0
		x"0A",x"E0",x"10",x"B0",x"F7",x"9D",x"93",x"02", -- 0x24C8
		x"E8",x"D0",x"F1",x"9D",x"93",x"02",x"20",x"94", -- 0x24D0
		x"E5",x"20",x"90",x"E7",x"8A",x"D0",x"CD",x"60", -- 0x24D8
		x"AD",x"A9",x"02",x"AC",x"AA",x"02",x"85",x"33", -- 0x24E0
		x"84",x"34",x"A0",x"00",x"20",x"C9",x"E6",x"AE", -- 0x24E8
		x"5B",x"02",x"D0",x"05",x"91",x"33",x"4C",x"05", -- 0x24F0
		x"E5",x"D1",x"33",x"F0",x"08",x"EE",x"5C",x"02", -- 0x24F8
		x"D0",x"03",x"EE",x"5D",x"02",x"20",x"6C",x"E5", -- 0x2500
		x"90",x"E2",x"60",x"10",x"07",x"53",x"65",x"61", -- 0x2508
		x"72",x"63",x"68",x"69",x"6E",x"67",x"20",x"2E", -- 0x2510
		x"2E",x"00",x"10",x"07",x"4C",x"6F",x"61",x"64", -- 0x2518
		x"69",x"6E",x"67",x"20",x"2E",x"2E",x"00",x"0A", -- 0x2520
		x"0D",x"45",x"72",x"72",x"6F",x"72",x"73",x"20", -- 0x2528
		x"66",x"6F",x"75",x"6E",x"64",x"0D",x"0A",x"00", -- 0x2530
		x"10",x"07",x"46",x"6F",x"75",x"6E",x"64",x"20", -- 0x2538
		x"2E",x"2E",x"00",x"10",x"07",x"56",x"65",x"72", -- 0x2540
		x"69",x"66",x"79",x"69",x"6E",x"67",x"20",x"2E", -- 0x2548
		x"2E",x"00",x"20",x"56",x"65",x"72",x"69",x"66", -- 0x2550
		x"79",x"20",x"65",x"72",x"72",x"6F",x"72",x"73", -- 0x2558
		x"20",x"64",x"65",x"74",x"65",x"63",x"74",x"65", -- 0x2560
		x"64",x"0D",x"0A",x"00",x"A5",x"33",x"CD",x"AB", -- 0x2568
		x"02",x"A5",x"34",x"ED",x"AC",x"02",x"E6",x"33", -- 0x2570
		x"D0",x"02",x"E6",x"34",x"60",x"A9",x"0B",x"A0", -- 0x2578
		x"E5",x"20",x"EA",x"E5",x"60",x"A9",x"45",x"A0", -- 0x2580
		x"E6",x"20",x"EA",x"E5",x"A9",x"7F",x"A0",x"02", -- 0x2588
		x"20",x"B6",x"E5",x"60",x"A9",x"38",x"A0",x"E5", -- 0x2590
		x"4C",x"AB",x"E5",x"AD",x"5B",x"02",x"D0",x"07", -- 0x2598
		x"A9",x"1A",x"A0",x"E5",x"4C",x"AB",x"E5",x"A9", -- 0x25A0
		x"43",x"A0",x"E5",x"20",x"EA",x"E5",x"A9",x"93", -- 0x25A8
		x"A0",x"02",x"20",x"B6",x"E5",x"60",x"20",x"65", -- 0x25B0
		x"F8",x"E8",x"A0",x"00",x"8C",x"5F",x"02",x"AD", -- 0x25B8
		x"AE",x"02",x"F0",x"13",x"C8",x"2C",x"AE",x"02", -- 0x25C0
		x"30",x"0D",x"C8",x"2C",x"AF",x"02",x"30",x"07", -- 0x25C8
		x"C8",x"2C",x"B0",x"02",x"30",x"01",x"C8",x"B9", -- 0x25D0
		x"E5",x"E5",x"8D",x"5E",x"02",x"A9",x"5E",x"A0", -- 0x25D8
		x"02",x"20",x"65",x"F8",x"60",x"42",x"43",x"53", -- 0x25E0
		x"49",x"52",x"20",x"F5",x"E5",x"A2",x"00",x"20", -- 0x25E8
		x"65",x"F8",x"E8",x"E8",x"60",x"48",x"AD",x"1F", -- 0x25F0
		x"02",x"D0",x"0A",x"A2",x"22",x"A9",x"10",x"9D", -- 0x25F8
		x"80",x"BB",x"CA",x"10",x"FA",x"68",x"60",x"20", -- 0x2600
		x"5A",x"E7",x"A9",x"24",x"20",x"5E",x"E6",x"A2", -- 0x2608
		x"09",x"BD",x"A7",x"02",x"20",x"5E",x"E6",x"CA", -- 0x2610
		x"D0",x"F7",x"BD",x"7F",x"02",x"F0",x"06",x"20", -- 0x2618
		x"5E",x"E6",x"E8",x"D0",x"F5",x"20",x"5E",x"E6", -- 0x2620
		x"A2",x"00",x"CA",x"D0",x"FD",x"60",x"AD",x"A9", -- 0x2628
		x"02",x"AC",x"AA",x"02",x"85",x"33",x"84",x"34", -- 0x2630
		x"A0",x"00",x"B1",x"33",x"20",x"5E",x"E6",x"20", -- 0x2638
		x"6C",x"E5",x"90",x"F6",x"60",x"10",x"07",x"53", -- 0x2640
		x"61",x"76",x"69",x"6E",x"67",x"20",x"2E",x"2E", -- 0x2648
		x"00",x"AD",x"B1",x"02",x"F0",x"07",x"A9",x"27", -- 0x2650
		x"A0",x"E5",x"20",x"B0",x"CC",x"60",x"85",x"2F", -- 0x2658
		x"8A",x"48",x"98",x"48",x"20",x"C0",x"E6",x"18", -- 0x2660
		x"A0",x"09",x"A9",x"00",x"F0",x"06",x"46",x"2F", -- 0x2668
		x"08",x"69",x"00",x"28",x"20",x"8B",x"E6",x"88", -- 0x2670
		x"D0",x"F4",x"49",x"01",x"4A",x"A0",x"04",x"20", -- 0x2678
		x"8B",x"E6",x"38",x"88",x"D0",x"F9",x"68",x"A8", -- 0x2680
		x"68",x"AA",x"60",x"48",x"08",x"AD",x"4D",x"02", -- 0x2688
		x"D0",x"0A",x"38",x"20",x"B2",x"E6",x"28",x"20", -- 0x2690
		x"B2",x"E6",x"68",x"60",x"20",x"B2",x"E6",x"A2", -- 0x2698
		x"0F",x"28",x"B0",x"02",x"A2",x"07",x"20",x"AB", -- 0x26A0
		x"E6",x"68",x"60",x"20",x"C0",x"E6",x"CA",x"D0", -- 0x26A8
		x"FA",x"60",x"A9",x"D0",x"A2",x"00",x"B0",x"02", -- 0x26B0
		x"0A",x"E8",x"8D",x"06",x"03",x"8E",x"07",x"03", -- 0x26B8
		x"AD",x"04",x"03",x"2C",x"0D",x"03",x"50",x"FB", -- 0x26C0
		x"60",x"98",x"48",x"8A",x"48",x"20",x"1C",x"E7", -- 0x26C8
		x"20",x"1C",x"E7",x"B0",x"FB",x"20",x"FF",x"E6", -- 0x26D0
		x"B0",x"16",x"A9",x"00",x"A0",x"08",x"20",x"FC", -- 0x26D8
		x"E6",x"08",x"66",x"2F",x"28",x"69",x"00",x"88", -- 0x26E0
		x"D0",x"F4",x"20",x"FC",x"E6",x"E9",x"00",x"4A", -- 0x26E8
		x"90",x"03",x"2E",x"B1",x"02",x"68",x"AA",x"68", -- 0x26F0
		x"A8",x"A5",x"2F",x"60",x"20",x"1C",x"E7",x"48", -- 0x26F8
		x"AD",x"4D",x"02",x"F0",x"15",x"20",x"1C",x"E7", -- 0x2700
		x"A2",x"02",x"90",x"02",x"A2",x"06",x"A9",x"00", -- 0x2708
		x"20",x"1C",x"E7",x"69",x"00",x"CA",x"D0",x"F8", -- 0x2710
		x"C9",x"04",x"68",x"60",x"48",x"AD",x"00",x"03", -- 0x2718
		x"AD",x"0D",x"03",x"29",x"10",x"F0",x"F9",x"AD", -- 0x2720
		x"09",x"03",x"48",x"A9",x"FF",x"8D",x"09",x"03", -- 0x2728
		x"68",x"C9",x"FE",x"68",x"60",x"20",x"FC",x"E6", -- 0x2730
		x"66",x"2F",x"A9",x"16",x"C5",x"2F",x"D0",x"F5", -- 0x2738
		x"AD",x"4D",x"02",x"F0",x"08",x"20",x"1C",x"E7", -- 0x2740
		x"20",x"1C",x"E7",x"B0",x"FB",x"A2",x"03",x"20", -- 0x2748
		x"C9",x"E6",x"C9",x"16",x"D0",x"DF",x"CA",x"D0", -- 0x2750
		x"F6",x"60",x"A2",x"02",x"A0",x"03",x"A9",x"16", -- 0x2758
		x"20",x"5E",x"E6",x"88",x"D0",x"F8",x"CA",x"D0", -- 0x2760
		x"F5",x"60",x"20",x"1A",x"EE",x"A0",x"06",x"78", -- 0x2768
		x"BE",x"82",x"E7",x"B9",x"89",x"E7",x"9D",x"00", -- 0x2770
		x"03",x"88",x"10",x"F4",x"A9",x"40",x"8D",x"00", -- 0x2778
		x"03",x"60",x"05",x"04",x"0B",x"02",x"0C",x"08", -- 0x2780
		x"0E",x"00",x"D0",x"C0",x"FF",x"10",x"F4",x"7F", -- 0x2788
		x"A0",x"00",x"A2",x"00",x"AD",x"7F",x"02",x"F0", -- 0x2790
		x"15",x"B9",x"7F",x"02",x"D9",x"93",x"02",x"F0", -- 0x2798
		x"01",x"E8",x"99",x"93",x"02",x"C8",x"C0",x"11", -- 0x27A0
		x"B0",x"04",x"48",x"68",x"D0",x"EB",x"60",x"4C", -- 0x27A8
		x"70",x"D0",x"A9",x"00",x"8D",x"4D",x"02",x"8D", -- 0x27B0
		x"AD",x"02",x"8D",x"AE",x"02",x"8D",x"5B",x"02", -- 0x27B8
		x"8D",x"5A",x"02",x"8D",x"5C",x"02",x"8D",x"5D", -- 0x27C0
		x"02",x"8D",x"B1",x"02",x"20",x"17",x"CF",x"24", -- 0x27C8
		x"28",x"10",x"DC",x"20",x"D0",x"D7",x"AA",x"A0", -- 0x27D0
		x"00",x"E8",x"CA",x"F0",x"0A",x"B1",x"91",x"99", -- 0x27D8
		x"7F",x"02",x"C8",x"C0",x"10",x"D0",x"F3",x"A9", -- 0x27E0
		x"00",x"99",x"7F",x"02",x"20",x"E8",x"00",x"F0", -- 0x27E8
		x"61",x"C9",x"2C",x"D0",x"BA",x"20",x"E2",x"00", -- 0x27F0
		x"F0",x"58",x"C9",x"2C",x"F0",x"F7",x"C9",x"C7", -- 0x27F8
		x"D0",x"05",x"8D",x"AD",x"02",x"B0",x"EE",x"C9", -- 0x2800
		x"53",x"D0",x"05",x"8D",x"4D",x"02",x"B0",x"E5", -- 0x2808
		x"C9",x"56",x"D0",x"05",x"8D",x"5B",x"02",x"B0", -- 0x2810
		x"DC",x"C9",x"4A",x"D0",x"05",x"8D",x"5A",x"02", -- 0x2818
		x"B0",x"D3",x"C9",x"41",x"F0",x"04",x"C9",x"45", -- 0x2820
		x"D0",x"47",x"85",x"0E",x"20",x"E2",x"00",x"A2", -- 0x2828
		x"80",x"8E",x"AE",x"02",x"20",x"53",x"E8",x"A5", -- 0x2830
		x"33",x"A4",x"34",x"A6",x"0E",x"E0",x"41",x"D0", -- 0x2838
		x"08",x"8D",x"A9",x"02",x"8C",x"AA",x"02",x"B0", -- 0x2840
		x"A3",x"8D",x"AB",x"02",x"8C",x"AC",x"02",x"4C", -- 0x2848
		x"EC",x"E7",x"60",x"20",x"03",x"CF",x"20",x"22", -- 0x2850
		x"D9",x"18",x"60",x"08",x"20",x"B2",x"E7",x"AD", -- 0x2858
		x"AD",x"02",x"0D",x"AE",x"02",x"D0",x"0A",x"AD", -- 0x2860
		x"5A",x"02",x"F0",x"08",x"AD",x"5B",x"02",x"F0", -- 0x2868
		x"03",x"4C",x"70",x"D0",x"20",x"6A",x"E7",x"20", -- 0x2870
		x"7D",x"E5",x"20",x"AC",x"E4",x"2C",x"AE",x"02", -- 0x2878
		x"70",x"F8",x"AD",x"5A",x"02",x"F0",x"2C",x"AD", -- 0x2880
		x"AE",x"02",x"D0",x"EE",x"A5",x"9C",x"A4",x"9D", -- 0x2888
		x"38",x"E9",x"02",x"B0",x"01",x"88",x"8D",x"A9", -- 0x2890
		x"02",x"8C",x"AA",x"02",x"38",x"E5",x"9A",x"AA", -- 0x2898
		x"98",x"E5",x"9B",x"A8",x"18",x"8A",x"6D",x"AB", -- 0x28A0
		x"02",x"8D",x"AB",x"02",x"98",x"6D",x"AC",x"02", -- 0x28A8
		x"8D",x"AC",x"02",x"20",x"9B",x"E5",x"20",x"E0", -- 0x28B0
		x"E4",x"20",x"3D",x"E9",x"28",x"AD",x"5B",x"02", -- 0x28B8
		x"F0",x"11",x"AE",x"5C",x"02",x"AD",x"5D",x"02", -- 0x28C0
		x"20",x"C5",x"E0",x"A9",x"52",x"A0",x"E5",x"20", -- 0x28C8
		x"B0",x"CC",x"60",x"20",x"51",x"E6",x"AD",x"AE", -- 0x28D0
		x"02",x"F0",x"0E",x"AD",x"AD",x"02",x"F0",x"08", -- 0x28D8
		x"AD",x"B1",x"02",x"EA",x"EA",x"6C",x"A9",x"02", -- 0x28E0
		x"60",x"AE",x"AB",x"02",x"AD",x"AC",x"02",x"86", -- 0x28E8
		x"9C",x"85",x"9D",x"20",x"5F",x"C5",x"AD",x"AD", -- 0x28F0
		x"02",x"F0",x"08",x"AD",x"B1",x"02",x"EA",x"EA", -- 0x28F8
		x"4C",x"08",x"C7",x"20",x"08",x"C7",x"4C",x"A8", -- 0x2900
		x"C4",x"A5",x"9A",x"A4",x"9B",x"8D",x"A9",x"02", -- 0x2908
		x"8C",x"AA",x"02",x"A5",x"9C",x"A4",x"9D",x"8D", -- 0x2910
		x"AB",x"02",x"8C",x"AC",x"02",x"08",x"20",x"B2", -- 0x2918
		x"E7",x"AD",x"5A",x"02",x"0D",x"5B",x"02",x"F0", -- 0x2920
		x"03",x"4C",x"70",x"D0",x"20",x"6A",x"E7",x"20", -- 0x2928
		x"85",x"E5",x"20",x"07",x"E6",x"20",x"2E",x"E6", -- 0x2930
		x"20",x"3D",x"E9",x"28",x"60",x"20",x"F5",x"E5", -- 0x2938
		x"20",x"AA",x"F9",x"4C",x"E0",x"ED",x"20",x"53", -- 0x2940
		x"E8",x"6C",x"33",x"00",x"A2",x"00",x"86",x"0C", -- 0x2948
		x"86",x"0D",x"F0",x"13",x"A2",x"03",x"0A",x"0A", -- 0x2950
		x"0A",x"0A",x"0A",x"26",x"0C",x"26",x"0D",x"90", -- 0x2958
		x"03",x"4C",x"39",x"DC",x"CA",x"10",x"F3",x"20", -- 0x2960
		x"E2",x"00",x"C9",x"80",x"B0",x"0E",x"09",x"80", -- 0x2968
		x"49",x"B0",x"C9",x"0A",x"90",x"DE",x"69",x"88", -- 0x2970
		x"C9",x"FA",x"B0",x"D8",x"A5",x"0D",x"A4",x"0C", -- 0x2978
		x"60",x"20",x"4C",x"E9",x"4C",x"40",x"DF",x"08", -- 0x2980
		x"20",x"57",x"EA",x"A9",x"40",x"8D",x"AE",x"02", -- 0x2988
		x"A5",x"28",x"8D",x"AF",x"02",x"A5",x"29",x"8D", -- 0x2990
		x"B0",x"02",x"20",x"85",x"E5",x"20",x"07",x"E6", -- 0x2998
		x"20",x"9E",x"EA",x"20",x"2E",x"E6",x"24",x"28", -- 0x29A0
		x"10",x"22",x"A0",x"00",x"B1",x"0C",x"F0",x"17", -- 0x29A8
		x"AA",x"A0",x"02",x"B1",x"0C",x"99",x"D0",x"00", -- 0x29B0
		x"88",x"D0",x"F8",x"E8",x"CA",x"F0",x"08",x"B1", -- 0x29B8
		x"D1",x"20",x"5E",x"E6",x"C8",x"D0",x"F5",x"20", -- 0x29C0
		x"42",x"EA",x"90",x"DE",x"20",x"3D",x"E9",x"28", -- 0x29C8
		x"60",x"20",x"50",x"D6",x"08",x"20",x"57",x"EA", -- 0x29D0
		x"20",x"7D",x"E5",x"20",x"AC",x"E4",x"2C",x"AE", -- 0x29D8
		x"02",x"50",x"F8",x"AD",x"AF",x"02",x"45",x"28", -- 0x29E0
		x"D0",x"F1",x"AD",x"B0",x"02",x"45",x"29",x"D0", -- 0x29E8
		x"EA",x"20",x"9B",x"E5",x"A0",x"02",x"B1",x"CE", -- 0x29F0
		x"CD",x"A9",x"02",x"C8",x"B1",x"CE",x"ED",x"AA", -- 0x29F8
		x"02",x"B0",x"06",x"20",x"3D",x"E9",x"4C",x"7C", -- 0x2A00
		x"C4",x"20",x"9E",x"EA",x"20",x"E0",x"E4",x"24", -- 0x2A08
		x"28",x"10",x"27",x"A0",x"00",x"B1",x"0C",x"F0", -- 0x2A10
		x"1C",x"20",x"AB",x"D5",x"A0",x"00",x"AA",x"E8", -- 0x2A18
		x"CA",x"F0",x"08",x"20",x"C9",x"E6",x"91",x"D1", -- 0x2A20
		x"C8",x"D0",x"F5",x"A0",x"02",x"B9",x"D0",x"00", -- 0x2A28
		x"91",x"0C",x"88",x"D0",x"F8",x"20",x"42",x"EA", -- 0x2A30
		x"90",x"D9",x"20",x"3D",x"E9",x"20",x"51",x"E6", -- 0x2A38
		x"28",x"60",x"18",x"A9",x"03",x"65",x"0C",x"85", -- 0x2A40
		x"0C",x"90",x"02",x"E6",x"0D",x"A8",x"A5",x"0D", -- 0x2A48
		x"CC",x"AB",x"02",x"ED",x"AC",x"02",x"60",x"A9", -- 0x2A50
		x"40",x"85",x"2B",x"20",x"88",x"D1",x"A9",x"00", -- 0x2A58
		x"85",x"2B",x"A0",x"03",x"B1",x"CE",x"8D",x"AA", -- 0x2A60
		x"02",x"88",x"B1",x"CE",x"8D",x"A9",x"02",x"D0", -- 0x2A68
		x"03",x"CE",x"AA",x"02",x"CE",x"A9",x"02",x"20", -- 0x2A70
		x"65",x"D0",x"A5",x"29",x"48",x"A5",x"28",x"48", -- 0x2A78
		x"20",x"B2",x"E7",x"68",x"85",x"28",x"68",x"85", -- 0x2A80
		x"29",x"AD",x"5B",x"02",x"0D",x"AD",x"02",x"0D", -- 0x2A88
		x"AE",x"02",x"0D",x"5A",x"02",x"F0",x"03",x"4C", -- 0x2A90
		x"70",x"D0",x"20",x"6A",x"E7",x"60",x"18",x"A5", -- 0x2A98
		x"CE",x"6D",x"A9",x"02",x"8D",x"AB",x"02",x"A5", -- 0x2AA0
		x"CF",x"6D",x"AA",x"02",x"8D",x"AC",x"02",x"A0", -- 0x2AA8
		x"04",x"B1",x"CE",x"20",x"88",x"D2",x"8D",x"A9", -- 0x2AB0
		x"02",x"8C",x"AA",x"02",x"85",x"0C",x"84",x"0D", -- 0x2AB8
		x"60",x"3F",x"FB",x"17",x"FC",x"CF",x"FB",x"C7", -- 0x2AC0
		x"F0",x"FC",x"F0",x"0F",x"F1",x"7E",x"F3",x"1C", -- 0x2AC8
		x"F1",x"67",x"F2",x"2C",x"F1",x"03",x"F2",x"0F", -- 0x2AD0
		x"F2",x"03",x"04",x"04",x"03",x"03",x"03",x"02", -- 0x2AD8
		x"01",x"03",x"03",x"01",x"01",x"00",x"00",x"00", -- 0x2AE0
		x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x2AE8
		x"AD",x"C0",x"02",x"29",x"01",x"D0",x"05",x"A2", -- 0x2AF0
		x"A3",x"4C",x"7E",x"C4",x"C0",x"4E",x"B0",x"03", -- 0x2AF8
		x"4C",x"70",x"D0",x"C0",x"66",x"B0",x"F9",x"98", -- 0x2B00
		x"38",x"E9",x"4E",x"A8",x"B9",x"C2",x"EA",x"48", -- 0x2B08
		x"B9",x"C1",x"EA",x"48",x"98",x"4A",x"A8",x"B9", -- 0x2B10
		x"D9",x"EA",x"48",x"B9",x"E5",x"EA",x"8D",x"C3", -- 0x2B18
		x"02",x"A9",x"00",x"8D",x"F0",x"02",x"20",x"03", -- 0x2B20
		x"CF",x"AD",x"C3",x"02",x"D0",x"06",x"20",x"22", -- 0x2B28
		x"D9",x"4C",x"3B",x"EB",x"A5",x"D0",x"C9",x"90", -- 0x2B30
		x"20",x"2A",x"D9",x"AC",x"F0",x"02",x"A5",x"33", -- 0x2B38
		x"99",x"E1",x"02",x"A5",x"34",x"99",x"E2",x"02", -- 0x2B40
		x"C8",x"C8",x"8C",x"F0",x"02",x"68",x"A8",x"88", -- 0x2B48
		x"F0",x"08",x"98",x"48",x"20",x"65",x"D0",x"4C", -- 0x2B50
		x"26",x"EB",x"A9",x"00",x"8D",x"E0",x"02",x"68", -- 0x2B58
		x"AA",x"68",x"A8",x"A9",x"EB",x"48",x"A9",x"6D", -- 0x2B60
		x"48",x"98",x"48",x"8A",x"48",x"60",x"A9",x"01", -- 0x2B68
		x"2C",x"E0",x"02",x"F0",x"F8",x"4C",x"36",x"D3", -- 0x2B70
		x"AD",x"DF",x"02",x"10",x"0B",x"08",x"29",x"7F", -- 0x2B78
		x"48",x"A9",x"00",x"8D",x"DF",x"02",x"68",x"28", -- 0x2B80
		x"60",x"C4",x"9D",x"B0",x"02",x"38",x"60",x"D0", -- 0x2B88
		x"06",x"C5",x"9C",x"90",x"F9",x"F0",x"F7",x"20", -- 0x2B90
		x"B5",x"EB",x"90",x"F2",x"AA",x"AD",x"C0",x"02", -- 0x2B98
		x"29",x"02",x"08",x"8A",x"28",x"D0",x"E6",x"98", -- 0x2BA0
		x"48",x"38",x"E9",x"1C",x"A8",x"8A",x"20",x"B5", -- 0x2BA8
		x"EB",x"68",x"A8",x"8A",x"60",x"CC",x"C2",x"02", -- 0x2BB0
		x"90",x"02",x"F0",x"01",x"60",x"CD",x"C1",x"02", -- 0x2BB8
		x"60",x"AC",x"C2",x"02",x"AD",x"C1",x"02",x"D0", -- 0x2BC0
		x"01",x"88",x"38",x"E9",x"01",x"60",x"20",x"03", -- 0x2BC8
		x"CF",x"20",x"22",x"D9",x"A5",x"33",x"A4",x"34", -- 0x2BD0
		x"20",x"89",x"EB",x"90",x"03",x"4C",x"7C",x"C4", -- 0x2BD8
		x"85",x"A6",x"84",x"A7",x"4C",x"0F",x"C7",x"AD", -- 0x2BE0
		x"60",x"02",x"D0",x"F1",x"AD",x"C0",x"02",x"48", -- 0x2BE8
		x"29",x"01",x"F0",x"05",x"A2",x"A3",x"4C",x"7E", -- 0x2BF0
		x"C4",x"68",x"29",x"FD",x"8D",x"C0",x"02",x"20", -- 0x2BF8
		x"C1",x"EB",x"48",x"98",x"18",x"69",x"1C",x"A8", -- 0x2C00
		x"68",x"4C",x"E0",x"EB",x"20",x"C1",x"EB",x"20", -- 0x2C08
		x"89",x"EB",x"B0",x"C9",x"48",x"AD",x"C0",x"02", -- 0x2C10
		x"09",x"02",x"8D",x"C0",x"02",x"68",x"4C",x"E0", -- 0x2C18
		x"EB",x"AD",x"C0",x"02",x"A8",x"29",x"01",x"F0", -- 0x2C20
		x"09",x"98",x"29",x"FE",x"8D",x"C0",x"02",x"20", -- 0x2C28
		x"67",x"F9",x"60",x"AD",x"C0",x"02",x"48",x"29", -- 0x2C30
		x"02",x"F0",x"B9",x"68",x"09",x"01",x"8D",x"C0", -- 0x2C38
		x"02",x"20",x"20",x"F9",x"60",x"20",x"62",x"D0", -- 0x2C40
		x"20",x"17",x"CF",x"A5",x"34",x"48",x"A5",x"33", -- 0x2C48
		x"48",x"20",x"22",x"D9",x"A5",x"33",x"8D",x"E1", -- 0x2C50
		x"02",x"A5",x"34",x"8D",x"E2",x"02",x"68",x"85", -- 0x2C58
		x"33",x"68",x"85",x"34",x"20",x"65",x"D0",x"20", -- 0x2C60
		x"17",x"CF",x"A5",x"34",x"48",x"A5",x"33",x"48", -- 0x2C68
		x"20",x"22",x"D9",x"A5",x"34",x"8D",x"E4",x"02", -- 0x2C70
		x"A5",x"33",x"8D",x"E3",x"02",x"68",x"85",x"33", -- 0x2C78
		x"68",x"85",x"34",x"20",x"C8",x"F1",x"AC",x"E1", -- 0x2C80
		x"02",x"AD",x"E0",x"02",x"29",x"01",x"D0",x"09", -- 0x2C88
		x"AD",x"E2",x"02",x"20",x"99",x"D4",x"4C",x"5F", -- 0x2C90
		x"D0",x"4C",x"C2",x"D8",x"E6",x"E9",x"D0",x"02", -- 0x2C98
		x"E6",x"EA",x"AD",x"60",x"EA",x"C9",x"20",x"F0", -- 0x2CA0
		x"F3",x"20",x"B9",x"EC",x"60",x"2C",x"60",x"EA", -- 0x2CA8
		x"2C",x"60",x"EA",x"60",x"80",x"4F",x"C7",x"52", -- 0x2CB0
		x"58",x"C9",x"C8",x"F0",x"0E",x"C9",x"27",x"F0", -- 0x2CB8
		x"0A",x"C9",x"3A",x"B0",x"06",x"38",x"E9",x"30", -- 0x2CC0
		x"38",x"E9",x"D0",x"60",x"D8",x"A2",x"FF",x"86", -- 0x2CC8
		x"A9",x"9A",x"A9",x"CC",x"A0",x"EC",x"85",x"1B", -- 0x2CD0
		x"84",x"1C",x"A9",x"4C",x"85",x"1A",x"85",x"C3", -- 0x2CD8
		x"85",x"21",x"8D",x"FB",x"02",x"A9",x"36",x"A0", -- 0x2CE0
		x"D3",x"85",x"22",x"84",x"23",x"8D",x"FC",x"02", -- 0x2CE8
		x"8C",x"FD",x"02",x"8D",x"F5",x"02",x"8C",x"F6", -- 0x2CF0
		x"02",x"A2",x"1C",x"BD",x"9B",x"EC",x"95",x"E1", -- 0x2CF8
		x"CA",x"D0",x"F8",x"A9",x"03",x"85",x"C2",x"8A", -- 0x2D00
		x"85",x"D7",x"85",x"87",x"85",x"2F",x"48",x"85", -- 0x2D08
		x"2E",x"8D",x"F2",x"02",x"A2",x"88",x"86",x"85", -- 0x2D10
		x"A8",x"A9",x"02",x"8D",x"C0",x"02",x"A9",x"28", -- 0x2D18
		x"8D",x"57",x"02",x"A9",x"50",x"8D",x"56",x"02", -- 0x2D20
		x"A9",x"00",x"85",x"30",x"8D",x"58",x"02",x"8D", -- 0x2D28
		x"59",x"02",x"20",x"3E",x"C8",x"20",x"CE",x"CC", -- 0x2D30
		x"A9",x"96",x"A0",x"ED",x"20",x"B0",x"CC",x"20", -- 0x2D38
		x"F0",x"CB",x"A2",x"00",x"A0",x"05",x"86",x"9A", -- 0x2D40
		x"84",x"9B",x"A0",x"00",x"98",x"91",x"9A",x"E6", -- 0x2D48
		x"9A",x"D0",x"02",x"E6",x"9B",x"20",x"F0",x"C6", -- 0x2D50
		x"A5",x"9A",x"A4",x"9B",x"20",x"44",x"C4",x"20", -- 0x2D58
		x"F0",x"CB",x"A5",x"A6",x"38",x"E5",x"9A",x"AA", -- 0x2D60
		x"A5",x"A7",x"E5",x"9B",x"20",x"C5",x"E0",x"A9", -- 0x2D68
		x"88",x"A0",x"ED",x"20",x"B0",x"CC",x"A9",x"B0", -- 0x2D70
		x"A0",x"CC",x"85",x"1B",x"84",x"1C",x"A9",x"10", -- 0x2D78
		x"8D",x"F8",x"02",x"4C",x"A8",x"C4",x"00",x"00", -- 0x2D80
		x"20",x"42",x"59",x"54",x"45",x"53",x"20",x"46", -- 0x2D88
		x"52",x"45",x"45",x"0A",x"0D",x"00",x"4F",x"52", -- 0x2D90
		x"49",x"43",x"20",x"45",x"58",x"54",x"45",x"4E", -- 0x2D98
		x"44",x"45",x"44",x"20",x"42",x"41",x"53",x"49", -- 0x2DA0
		x"43",x"20",x"56",x"31",x"2E",x"31",x"0D",x"0A", -- 0x2DA8
		x"60",x"20",x"31",x"39",x"38",x"33",x"20",x"54", -- 0x2DB0
		x"41",x"4E",x"47",x"45",x"52",x"49",x"4E",x"45", -- 0x2DB8
		x"0D",x"0A",x"00",x"00",x"A2",x"00",x"A0",x"00", -- 0x2DC0
		x"C4",x"10",x"D0",x"04",x"E4",x"11",x"F0",x"0F", -- 0x2DC8
		x"B1",x"0C",x"91",x"0E",x"C8",x"D0",x"F1",x"E6", -- 0x2DD0
		x"0D",x"E6",x"0F",x"E8",x"4C",x"C8",x"ED",x"60", -- 0x2DD8
		x"48",x"20",x"8C",x"EE",x"A9",x"00",x"A2",x"00", -- 0x2DE0
		x"A0",x"03",x"20",x"AB",x"EE",x"A9",x"01",x"A0", -- 0x2DE8
		x"19",x"20",x"AB",x"EE",x"A9",x"00",x"8D",x"71", -- 0x2DF0
		x"02",x"AD",x"0B",x"03",x"29",x"7F",x"09",x"40", -- 0x2DF8
		x"8D",x"0B",x"03",x"A9",x"C0",x"8D",x"0E",x"03", -- 0x2E00
		x"A9",x"10",x"8D",x"06",x"03",x"8D",x"04",x"03", -- 0x2E08
		x"A9",x"27",x"8D",x"07",x"03",x"8D",x"05",x"03", -- 0x2E10
		x"68",x"60",x"48",x"A9",x"40",x"8D",x"0E",x"03", -- 0x2E18
		x"68",x"60",x"48",x"AD",x"0D",x"03",x"29",x"40", -- 0x2E20
		x"F0",x"06",x"8D",x"0D",x"03",x"20",x"34",x"EE", -- 0x2E28
		x"68",x"4C",x"4A",x"02",x"48",x"8A",x"48",x"98", -- 0x2E30
		x"48",x"A0",x"00",x"B9",x"72",x"02",x"38",x"E9", -- 0x2E38
		x"01",x"99",x"72",x"02",x"C8",x"B9",x"72",x"02", -- 0x2E40
		x"E9",x"00",x"99",x"72",x"02",x"C8",x"C0",x"06", -- 0x2E48
		x"D0",x"E9",x"A9",x"00",x"20",x"9D",x"EE",x"C0", -- 0x2E50
		x"00",x"D0",x"10",x"A2",x"00",x"A0",x"03",x"20", -- 0x2E58
		x"AB",x"EE",x"20",x"95",x"F4",x"8A",x"10",x"03", -- 0x2E60
		x"8E",x"DF",x"02",x"A9",x"01",x"20",x"9D",x"EE", -- 0x2E68
		x"C0",x"00",x"D0",x"12",x"A2",x"00",x"A0",x"19", -- 0x2E70
		x"20",x"AB",x"EE",x"AD",x"71",x"02",x"49",x"01", -- 0x2E78
		x"8D",x"71",x"02",x"20",x"01",x"F8",x"68",x"A8", -- 0x2E80
		x"68",x"AA",x"68",x"60",x"48",x"98",x"48",x"A0", -- 0x2E88
		x"05",x"A9",x"00",x"99",x"72",x"02",x"88",x"10", -- 0x2E90
		x"FA",x"68",x"A8",x"68",x"60",x"48",x"0A",x"A8", -- 0x2E98
		x"78",x"B9",x"72",x"02",x"BE",x"73",x"02",x"58", -- 0x2EA0
		x"A8",x"68",x"60",x"48",x"8A",x"48",x"98",x"48", -- 0x2EA8
		x"BA",x"BD",x"03",x"01",x"0A",x"A8",x"68",x"48", -- 0x2EB0
		x"78",x"99",x"72",x"02",x"BD",x"02",x"01",x"99", -- 0x2EB8
		x"73",x"02",x"58",x"68",x"A8",x"68",x"AA",x"68", -- 0x2EC0
		x"60",x"20",x"AB",x"EE",x"20",x"9D",x"EE",x"C0", -- 0x2EC8
		x"00",x"D0",x"F9",x"E0",x"00",x"D0",x"F5",x"60", -- 0x2ED0
		x"AD",x"13",x"02",x"8D",x"14",x"02",x"4E",x"12", -- 0x2ED8
		x"02",x"6E",x"12",x"02",x"6E",x"12",x"02",x"60", -- 0x2EE0
		x"48",x"98",x"48",x"20",x"DE",x"EE",x"20",x"49", -- 0x2EE8
		x"F0",x"20",x"24",x"F0",x"68",x"A8",x"68",x"60", -- 0x2EF0
		x"D8",x"20",x"D8",x"EE",x"2C",x"E2",x"02",x"10", -- 0x2EF8
		x"0A",x"A9",x"FF",x"4D",x"E1",x"02",x"AA",x"E8", -- 0x2F00
		x"8E",x"E1",x"02",x"2C",x"E4",x"02",x"10",x"0A", -- 0x2F08
		x"A9",x"FF",x"4D",x"E3",x"02",x"AA",x"E8",x"8E", -- 0x2F10
		x"E3",x"02",x"AD",x"E1",x"02",x"CD",x"E3",x"02", -- 0x2F18
		x"90",x"0F",x"AE",x"E1",x"02",x"F0",x"09",x"AD", -- 0x2F20
		x"E3",x"02",x"20",x"40",x"EF",x"20",x"84",x"EF", -- 0x2F28
		x"60",x"AE",x"E3",x"02",x"F0",x"09",x"AD",x"E1", -- 0x2F30
		x"02",x"20",x"40",x"EF",x"20",x"5C",x"EF",x"60", -- 0x2F38
		x"85",x"0D",x"8E",x"00",x"02",x"A9",x"00",x"85", -- 0x2F40
		x"0C",x"8D",x"01",x"02",x"20",x"C8",x"EF",x"20", -- 0x2F48
		x"FA",x"EF",x"A9",x"00",x"85",x"0E",x"85",x"0F", -- 0x2F50
		x"8D",x"00",x"02",x"60",x"2C",x"E4",x"02",x"10", -- 0x2F58
		x"06",x"20",x"95",x"F0",x"4C",x"6A",x"EF",x"20", -- 0x2F60
		x"89",x"F0",x"20",x"AC",x"EF",x"F0",x"0E",x"2C", -- 0x2F68
		x"E2",x"02",x"10",x"06",x"20",x"B2",x"F0",x"4C", -- 0x2F70
		x"7D",x"EF",x"20",x"A1",x"F0",x"20",x"16",x"F0", -- 0x2F78
		x"CA",x"D0",x"D9",x"60",x"2C",x"E2",x"02",x"10", -- 0x2F80
		x"06",x"20",x"B2",x"F0",x"4C",x"92",x"EF",x"20", -- 0x2F88
		x"A1",x"F0",x"20",x"AC",x"EF",x"F0",x"0E",x"2C", -- 0x2F90
		x"E4",x"02",x"10",x"06",x"20",x"95",x"F0",x"4C", -- 0x2F98
		x"A5",x"EF",x"20",x"89",x"F0",x"20",x"16",x"F0", -- 0x2FA0
		x"CA",x"D0",x"D9",x"60",x"D8",x"18",x"A5",x"0E", -- 0x2FA8
		x"65",x"0C",x"85",x"0E",x"A5",x"0F",x"65",x"0D", -- 0x2FB0
		x"85",x"0F",x"24",x"0E",x"10",x"03",x"18",x"69", -- 0x2FB8
		x"01",x"CD",x"00",x"02",x"8D",x"00",x"02",x"60", -- 0x2FC0
		x"48",x"8A",x"48",x"98",x"48",x"A9",x"00",x"85", -- 0x2FC8
		x"0E",x"85",x"0F",x"A2",x"10",x"06",x"0C",x"26", -- 0x2FD0
		x"0D",x"26",x"0E",x"26",x"0F",x"A5",x"0E",x"38", -- 0x2FD8
		x"ED",x"00",x"02",x"A8",x"A5",x"0F",x"ED",x"01", -- 0x2FE0
		x"02",x"90",x"06",x"E6",x"0C",x"84",x"0E",x"85", -- 0x2FE8
		x"0F",x"CA",x"D0",x"E1",x"68",x"A8",x"68",x"AA", -- 0x2FF0
		x"68",x"60",x"48",x"0E",x"00",x"02",x"2E",x"01", -- 0x2FF8
		x"02",x"AD",x"00",x"02",x"38",x"E5",x"0E",x"AD", -- 0x3000
		x"01",x"02",x"E5",x"0F",x"B0",x"06",x"E6",x"0C", -- 0x3008
		x"D0",x"02",x"E6",x"0D",x"68",x"60",x"2C",x"14", -- 0x3010
		x"02",x"18",x"10",x"04",x"20",x"24",x"F0",x"38", -- 0x3018
		x"2E",x"14",x"02",x"60",x"A0",x"00",x"B1",x"10", -- 0x3020
		x"29",x"40",x"F0",x"1C",x"AD",x"15",x"02",x"2C", -- 0x3028
		x"12",x"02",x"30",x"0E",x"70",x"07",x"49",x"FF", -- 0x3030
		x"31",x"10",x"91",x"10",x"60",x"11",x"10",x"91", -- 0x3038
		x"10",x"60",x"70",x"04",x"51",x"10",x"91",x"10", -- 0x3040
		x"60",x"D8",x"48",x"98",x"48",x"20",x"31",x"F7", -- 0x3048
		x"18",x"69",x"00",x"85",x"10",x"98",x"69",x"A0", -- 0x3050
		x"85",x"11",x"A9",x"00",x"85",x"0D",x"8D",x"01", -- 0x3058
		x"02",x"86",x"0C",x"A9",x"06",x"8D",x"00",x"02", -- 0x3060
		x"20",x"C8",x"EF",x"18",x"A5",x"0C",x"65",x"10", -- 0x3068
		x"85",x"10",x"A9",x"00",x"65",x"11",x"85",x"11", -- 0x3070
		x"A9",x"20",x"A4",x"0E",x"F0",x"04",x"4A",x"88", -- 0x3078
		x"90",x"FA",x"8D",x"15",x"02",x"68",x"A8",x"68", -- 0x3080
		x"60",x"18",x"A5",x"10",x"69",x"28",x"85",x"10", -- 0x3088
		x"90",x"02",x"E6",x"11",x"60",x"38",x"A5",x"10", -- 0x3090
		x"E9",x"28",x"85",x"10",x"B0",x"02",x"C6",x"11", -- 0x3098
		x"60",x"4E",x"15",x"02",x"90",x"0B",x"A9",x"20", -- 0x30A0
		x"8D",x"15",x"02",x"E6",x"10",x"D0",x"02",x"E6", -- 0x30A8
		x"11",x"60",x"0E",x"15",x"02",x"2C",x"15",x"02", -- 0x30B0
		x"50",x"0D",x"A9",x"01",x"8D",x"15",x"02",x"A5", -- 0x30B8
		x"10",x"D0",x"02",x"C6",x"11",x"C6",x"10",x"60", -- 0x30C0
		x"A9",x"04",x"A2",x"E5",x"20",x"F8",x"F2",x"B0", -- 0x30C8
		x"28",x"AD",x"E5",x"02",x"8D",x"12",x"02",x"A9", -- 0x30D0
		x"F0",x"A2",x"E1",x"20",x"F8",x"F2",x"B0",x"19", -- 0x30D8
		x"A9",x"C8",x"A2",x"E3",x"20",x"F8",x"F2",x"B0", -- 0x30E0
		x"10",x"AE",x"E1",x"02",x"8E",x"19",x"02",x"AC", -- 0x30E8
		x"E3",x"02",x"8C",x"1A",x"02",x"20",x"E8",x"EE", -- 0x30F0
		x"60",x"EE",x"E0",x"02",x"60",x"20",x"0A",x"F3", -- 0x30F8
		x"B0",x"0A",x"AE",x"19",x"02",x"AC",x"1A",x"02", -- 0x3100
		x"20",x"E8",x"EE",x"60",x"EE",x"E0",x"02",x"60", -- 0x3108
		x"20",x"0A",x"F3",x"B0",x"04",x"20",x"F8",x"EE", -- 0x3110
		x"60",x"EE",x"E0",x"02",x"60",x"AE",x"E2",x"02", -- 0x3118
		x"D0",x"07",x"AE",x"E1",x"02",x"8E",x"13",x"02", -- 0x3120
		x"60",x"EE",x"E0",x"02",x"60",x"AE",x"E2",x"02", -- 0x3128
		x"D0",x"3B",x"AE",x"E1",x"02",x"E0",x"20",x"90", -- 0x3130
		x"34",x"E0",x"80",x"B0",x"30",x"A9",x"02",x"A2", -- 0x3138
		x"E3",x"20",x"F8",x"F2",x"B0",x"27",x"A9",x"04", -- 0x3140
		x"A2",x"E5",x"20",x"F8",x"F2",x"B0",x"1E",x"AD", -- 0x3148
		x"19",x"02",x"C9",x"EB",x"B0",x"17",x"AD",x"1A", -- 0x3150
		x"02",x"C9",x"C1",x"B0",x"10",x"20",x"71",x"F1", -- 0x3158
		x"20",x"9B",x"F1",x"AE",x"19",x"02",x"AC",x"1A", -- 0x3160
		x"02",x"20",x"49",x"F0",x"60",x"EE",x"E0",x"02", -- 0x3168
		x"60",x"D8",x"AD",x"E5",x"02",x"8D",x"12",x"02", -- 0x3170
		x"20",x"DE",x"EE",x"AD",x"E1",x"02",x"85",x"0C", -- 0x3178
		x"A9",x"00",x"85",x"0D",x"A2",x"03",x"06",x"0C", -- 0x3180
		x"26",x"0D",x"CA",x"D0",x"F9",x"AD",x"E3",x"02", -- 0x3188
		x"0A",x"0A",x"18",x"69",x"98",x"18",x"65",x"0D", -- 0x3190
		x"85",x"0D",x"60",x"D8",x"A0",x"00",x"84",x"0F", -- 0x3198
		x"B1",x"0C",x"85",x"0E",x"20",x"5D",x"F3",x"26", -- 0x31A0
		x"0E",x"26",x"0E",x"A2",x"06",x"26",x"0E",x"90", -- 0x31A8
		x"03",x"20",x"24",x"F0",x"20",x"A1",x"F0",x"CA", -- 0x31B0
		x"D0",x"F3",x"20",x"6E",x"F3",x"20",x"89",x"F0", -- 0x31B8
		x"A4",x"0F",x"C8",x"C0",x"08",x"D0",x"D7",x"60", -- 0x31C0
		x"A9",x"F0",x"A2",x"E1",x"20",x"F8",x"F2",x"B0", -- 0x31C8
		x"2F",x"A9",x"C8",x"A2",x"E3",x"20",x"F8",x"F2", -- 0x31D0
		x"B0",x"26",x"AE",x"E1",x"02",x"8E",x"19",x"02", -- 0x31D8
		x"AC",x"E3",x"02",x"8C",x"1A",x"02",x"20",x"49", -- 0x31E0
		x"F0",x"A0",x"00",x"B1",x"10",x"2D",x"15",x"02", -- 0x31E8
		x"F0",x"05",x"A9",x"FF",x"4C",x"F9",x"F1",x"A9", -- 0x31F0
		x"00",x"8D",x"E1",x"02",x"8D",x"E2",x"02",x"60", -- 0x31F8
		x"EE",x"E0",x"02",x"60",x"A9",x"10",x"85",x"0C", -- 0x3200
		x"A9",x"00",x"85",x"0D",x"20",x"1C",x"F2",x"60", -- 0x3208
		x"A9",x"00",x"85",x"0C",x"A9",x"01",x"85",x"0D", -- 0x3210
		x"20",x"1C",x"F2",x"60",x"A9",x"08",x"A2",x"E1", -- 0x3218
		x"20",x"F8",x"F2",x"B0",x"3F",x"20",x"5D",x"F3", -- 0x3220
		x"AD",x"E1",x"02",x"05",x"0C",x"8D",x"02",x"02", -- 0x3228
		x"AE",x"1F",x"02",x"D0",x"12",x"A6",x"0D",x"9D", -- 0x3230
		x"6B",x"02",x"A9",x"A8",x"18",x"65",x"0D",x"AA", -- 0x3238
		x"A0",x"BB",x"A9",x"1B",x"4C",x"51",x"F2",x"A9", -- 0x3240
		x"00",x"18",x"65",x"0D",x"AA",x"A0",x"A0",x"A9", -- 0x3248
		x"C8",x"8D",x"00",x"02",x"86",x"10",x"84",x"11", -- 0x3250
		x"A9",x"01",x"8D",x"01",x"02",x"20",x"CD",x"F2", -- 0x3258
		x"20",x"6E",x"F3",x"60",x"EE",x"E0",x"02",x"60", -- 0x3260
		x"D8",x"AD",x"E3",x"02",x"8D",x"01",x"02",x"F0", -- 0x3268
		x"58",x"A0",x"00",x"AD",x"19",x"02",x"38",x"E9", -- 0x3270
		x"06",x"90",x"04",x"C8",x"4C",x"76",x"F2",x"98", -- 0x3278
		x"18",x"6D",x"E3",x"02",x"A8",x"AD",x"E4",x"02", -- 0x3280
		x"69",x"00",x"D0",x"3D",x"C0",x"29",x"B0",x"39", -- 0x3288
		x"AD",x"E6",x"02",x"D0",x"34",x"AD",x"E1",x"02", -- 0x3290
		x"8D",x"00",x"02",x"F0",x"2C",x"18",x"6D",x"1A", -- 0x3298
		x"02",x"A8",x"AD",x"E2",x"02",x"69",x"00",x"D0", -- 0x32A0
		x"20",x"C0",x"C9",x"B0",x"1C",x"C0",x"C8",x"D0", -- 0x32A8
		x"02",x"A0",x"00",x"8C",x"1A",x"02",x"AD",x"E5", -- 0x32B0
		x"02",x"8D",x"02",x"02",x"20",x"CD",x"F2",x"AC", -- 0x32B8
		x"1A",x"02",x"AE",x"19",x"02",x"20",x"49",x"F0", -- 0x32C0
		x"60",x"EE",x"E0",x"02",x"60",x"D8",x"AD",x"02", -- 0x32C8
		x"02",x"A0",x"00",x"91",x"10",x"C8",x"CC",x"01", -- 0x32D0
		x"02",x"D0",x"F8",x"20",x"89",x"F0",x"CE",x"00", -- 0x32D8
		x"02",x"D0",x"EB",x"60",x"8D",x"04",x"02",x"BD", -- 0x32E0
		x"01",x"02",x"D0",x"0A",x"BD",x"00",x"02",x"F0", -- 0x32E8
		x"05",x"CD",x"04",x"02",x"90",x"01",x"38",x"60", -- 0x32F0
		x"8D",x"04",x"02",x"BD",x"01",x"02",x"D0",x"08", -- 0x32F8
		x"BD",x"00",x"02",x"CD",x"04",x"02",x"90",x"01", -- 0x3300
		x"38",x"60",x"A9",x"04",x"A2",x"E5",x"20",x"F8", -- 0x3308
		x"F2",x"B0",x"49",x"18",x"AD",x"E1",x"02",x"6D", -- 0x3310
		x"19",x"02",x"8D",x"00",x"02",x"AD",x"E2",x"02", -- 0x3318
		x"69",x"00",x"8D",x"01",x"02",x"A2",x"00",x"A9", -- 0x3320
		x"F0",x"20",x"F8",x"F2",x"B0",x"2E",x"18",x"AD", -- 0x3328
		x"E3",x"02",x"6D",x"1A",x"02",x"8D",x"02",x"02", -- 0x3330
		x"AD",x"E4",x"02",x"69",x"00",x"8D",x"03",x"02", -- 0x3338
		x"A2",x"02",x"A9",x"C8",x"20",x"F8",x"F2",x"B0", -- 0x3340
		x"13",x"AD",x"E5",x"02",x"8D",x"12",x"02",x"AD", -- 0x3348
		x"00",x"02",x"8D",x"19",x"02",x"AD",x"02",x"02", -- 0x3350
		x"8D",x"1A",x"02",x"18",x"60",x"A5",x"10",x"8D", -- 0x3358
		x"16",x"02",x"A5",x"11",x"8D",x"17",x"02",x"AD", -- 0x3360
		x"15",x"02",x"8D",x"18",x"02",x"60",x"AD",x"16", -- 0x3368
		x"02",x"85",x"10",x"AD",x"17",x"02",x"85",x"11", -- 0x3370
		x"AD",x"18",x"02",x"8D",x"15",x"02",x"60",x"D8", -- 0x3378
		x"AD",x"E2",x"02",x"D0",x"3D",x"AD",x"E1",x"02", -- 0x3380
		x"F0",x"38",x"AD",x"19",x"02",x"CD",x"E1",x"02", -- 0x3388
		x"90",x"30",x"18",x"6D",x"E1",x"02",x"C9",x"F0", -- 0x3390
		x"B0",x"28",x"AD",x"1A",x"02",x"CD",x"E1",x"02", -- 0x3398
		x"90",x"20",x"18",x"6D",x"E1",x"02",x"C9",x"C8", -- 0x33A0
		x"B0",x"18",x"A2",x"E3",x"A9",x"04",x"20",x"F8", -- 0x33A8
		x"F2",x"B0",x"0F",x"AD",x"E3",x"02",x"8D",x"12", -- 0x33B0
		x"02",x"20",x"D8",x"EE",x"20",x"C6",x"F3",x"4C", -- 0x33B8
		x"C5",x"F3",x"EE",x"E0",x"02",x"60",x"20",x"5D", -- 0x33C0
		x"F3",x"AD",x"1A",x"02",x"38",x"ED",x"E1",x"02", -- 0x33C8
		x"A8",x"AE",x"19",x"02",x"20",x"49",x"F0",x"AD", -- 0x33D0
		x"E1",x"02",x"85",x"0F",x"20",x"85",x"F4",x"A9", -- 0x33D8
		x"80",x"8D",x"1B",x"02",x"8D",x"1D",x"02",x"A9", -- 0x33E0
		x"00",x"8D",x"1C",x"02",x"AD",x"E1",x"02",x"8D", -- 0x33E8
		x"1E",x"02",x"A9",x"00",x"85",x"0F",x"20",x"14", -- 0x33F0
		x"F4",x"20",x"44",x"F4",x"A5",x"0F",x"F0",x"03", -- 0x33F8
		x"20",x"16",x"F0",x"AD",x"1C",x"02",x"D0",x"EA", -- 0x3400
		x"AD",x"1E",x"02",x"CD",x"E1",x"02",x"D0",x"E2", -- 0x3408
		x"20",x"6E",x"F3",x"60",x"AD",x"1D",x"02",x"AE", -- 0x3410
		x"1E",x"02",x"20",x"74",x"F4",x"A5",x"0C",x"18", -- 0x3418
		x"6D",x"1B",x"02",x"8D",x"1B",x"02",x"AD",x"1C", -- 0x3420
		x"02",x"85",x"0C",x"65",x"0D",x"8D",x"1C",x"02", -- 0x3428
		x"C5",x"0C",x"F0",x"0F",x"B0",x"06",x"20",x"A1", -- 0x3430
		x"F0",x"4C",x"3F",x"F4",x"20",x"B2",x"F0",x"A9", -- 0x3438
		x"01",x"85",x"0F",x"60",x"AD",x"1B",x"02",x"AE", -- 0x3440
		x"1C",x"02",x"20",x"74",x"F4",x"38",x"AD",x"1D", -- 0x3448
		x"02",x"E5",x"0C",x"8D",x"1D",x"02",x"AD",x"1E", -- 0x3450
		x"02",x"85",x"0C",x"E5",x"0D",x"8D",x"1E",x"02", -- 0x3458
		x"C5",x"0C",x"F0",x"0F",x"B0",x"06",x"20",x"89", -- 0x3460
		x"F0",x"4C",x"6F",x"F4",x"20",x"95",x"F0",x"A9", -- 0x3468
		x"01",x"85",x"0F",x"60",x"85",x"0C",x"86",x"0D", -- 0x3470
		x"A6",x"0E",x"A5",x"0D",x"2A",x"66",x"0D",x"66", -- 0x3478
		x"0C",x"CA",x"D0",x"F6",x"60",x"E6",x"0F",x"A9", -- 0x3480
		x"00",x"85",x"0E",x"A9",x"01",x"0A",x"E6",x"0E", -- 0x3488
		x"C5",x"0F",x"90",x"F9",x"60",x"48",x"08",x"98", -- 0x3490
		x"48",x"D8",x"AD",x"08",x"02",x"10",x"1E",x"29", -- 0x3498
		x"87",x"8D",x"10",x"02",x"AE",x"0A",x"02",x"20", -- 0x34A0
		x"61",x"F5",x"CD",x"10",x"02",x"D0",x"0E",x"CE", -- 0x34A8
		x"0E",x"02",x"D0",x"33",x"AD",x"4F",x"02",x"8D", -- 0x34B0
		x"0E",x"02",x"4C",x"C6",x"F4",x"AD",x"4E",x"02", -- 0x34B8
		x"8D",x"0E",x"02",x"20",x"23",x"F5",x"20",x"EF", -- 0x34C0
		x"F4",x"AA",x"10",x"1D",x"48",x"AD",x"6A",x"02", -- 0x34C8
		x"29",x"08",x"D0",x"0F",x"68",x"48",x"C9",x"A0", -- 0x34D0
		x"90",x"06",x"20",x"14",x"FB",x"4C",x"E3",x"F4", -- 0x34D8
		x"20",x"2A",x"FB",x"68",x"4C",x"E9",x"F4",x"A9", -- 0x34E0
		x"00",x"AA",x"68",x"A8",x"28",x"68",x"60",x"AD", -- 0x34E8
		x"09",x"02",x"A8",x"A9",x"00",x"C0",x"A4",x"F0", -- 0x34F0
		x"04",x"C0",x"A7",x"D0",x"03",x"18",x"69",x"40", -- 0x34F8
		x"18",x"6D",x"08",x"02",x"10",x"1C",x"29",x"7F", -- 0x3500
		x"AA",x"BD",x"78",x"FF",x"2D",x"0C",x"02",x"10", -- 0x3508
		x"03",x"38",x"E9",x"20",x"29",x"7F",x"C0",x"A2", -- 0x3510
		x"D0",x"06",x"C9",x"40",x"30",x"02",x"29",x"1F", -- 0x3518
		x"09",x"80",x"60",x"A9",x"38",x"8D",x"0D",x"02", -- 0x3520
		x"8D",x"08",x"02",x"8D",x"09",x"02",x"A9",x"7F", -- 0x3528
		x"48",x"68",x"48",x"AA",x"A9",x"07",x"20",x"61", -- 0x3530
		x"F5",x"0D",x"0D",x"02",x"10",x"12",x"A2",x"00", -- 0x3538
		x"A0",x"20",x"CC",x"0D",x"02",x"D0",x"01",x"E8", -- 0x3540
		x"9D",x"08",x"02",x"68",x"48",x"9D",x"0A",x"02", -- 0x3548
		x"38",x"68",x"6A",x"48",x"38",x"AD",x"0D",x"02", -- 0x3550
		x"E9",x"08",x"8D",x"0D",x"02",x"10",x"D2",x"68", -- 0x3558
		x"60",x"48",x"A9",x"0E",x"20",x"90",x"F5",x"68", -- 0x3560
		x"29",x"07",x"AA",x"8D",x"11",x"02",x"09",x"B8", -- 0x3568
		x"8D",x"00",x"03",x"A0",x"04",x"88",x"D0",x"FD", -- 0x3570
		x"AD",x"00",x"03",x"29",x"08",x"D0",x"0D",x"CA", -- 0x3578
		x"8A",x"29",x"07",x"AA",x"CD",x"11",x"02",x"D0", -- 0x3580
		x"E5",x"A9",x"00",x"60",x"8A",x"09",x"80",x"60", -- 0x3588
		x"08",x"78",x"8D",x"0F",x"03",x"A8",x"8A",x"C0", -- 0x3590
		x"07",x"D0",x"02",x"09",x"40",x"48",x"AD",x"0C", -- 0x3598
		x"03",x"09",x"EE",x"8D",x"0C",x"03",x"29",x"11", -- 0x35A0
		x"09",x"CC",x"8D",x"0C",x"03",x"AA",x"68",x"8D", -- 0x35A8
		x"0F",x"03",x"8A",x"09",x"EC",x"8D",x"0C",x"03", -- 0x35B0
		x"29",x"11",x"09",x"CC",x"8D",x"0C",x"03",x"28", -- 0x35B8
		x"60",x"08",x"78",x"8D",x"01",x"03",x"AD",x"00", -- 0x35C0
		x"03",x"29",x"EF",x"8D",x"00",x"03",x"AD",x"00", -- 0x35C8
		x"03",x"09",x"10",x"8D",x"00",x"03",x"28",x"AD", -- 0x35D0
		x"0D",x"03",x"29",x"02",x"F0",x"F9",x"AD",x"0D", -- 0x35D8
		x"03",x"60",x"CF",x"CF",x"CF",x"CF",x"A3",x"CF", -- 0x35E0
		x"A6",x"CC",x"00",x"27",x"34",x"0F",x"66",x"99", -- 0x35E8
		x"60",x"CF",x"A7",x"B3",x"CF",x"A8",x"BE",x"CF", -- 0x35F0
		x"CF",x"CF",x"CF",x"CF",x"A5",x"A5",x"CF",x"A4", -- 0x35F8
		x"84",x"CF",x"29",x"1F",x"AA",x"BD",x"E2",x"F5", -- 0x3600
		x"18",x"69",x"2F",x"8D",x"61",x"02",x"A9",x"00", -- 0x3608
		x"69",x"F6",x"8D",x"62",x"02",x"AD",x"6A",x"02", -- 0x3610
		x"48",x"29",x"FE",x"8D",x"6A",x"02",x"68",x"29", -- 0x3618
		x"01",x"8D",x"51",x"02",x"A9",x"00",x"20",x"01", -- 0x3620
		x"F8",x"38",x"A9",x"00",x"6C",x"61",x"02",x"CE", -- 0x3628
		x"69",x"02",x"30",x"05",x"20",x"D7",x"F7",x"D0", -- 0x3630
		x"40",x"A9",x"27",x"8D",x"69",x"02",x"AD",x"68", -- 0x3638
		x"02",x"C9",x"01",x"F0",x"34",x"CE",x"68",x"02", -- 0x3640
		x"38",x"A5",x"12",x"E9",x"28",x"85",x"12",x"B0", -- 0x3648
		x"02",x"C6",x"13",x"4C",x"FE",x"F6",x"EE",x"69", -- 0x3650
		x"02",x"A2",x"27",x"EC",x"69",x"02",x"10",x"19", -- 0x3658
		x"20",x"0D",x"F7",x"AD",x"68",x"02",x"CD",x"7E", -- 0x3660
		x"02",x"F0",x"11",x"EE",x"68",x"02",x"18",x"A5", -- 0x3668
		x"12",x"69",x"28",x"85",x"12",x"90",x"02",x"E6", -- 0x3670
		x"13",x"4C",x"FE",x"F6",x"20",x"5D",x"F3",x"A2", -- 0x3678
		x"06",x"BD",x"77",x"02",x"95",x"0B",x"CA",x"D0", -- 0x3680
		x"F8",x"20",x"C4",x"ED",x"20",x"6E",x"F3",x"20", -- 0x3688
		x"1A",x"F7",x"4C",x"FE",x"F6",x"AE",x"7E",x"02", -- 0x3690
		x"AD",x"7A",x"02",x"85",x"12",x"AD",x"7B",x"02", -- 0x3698
		x"85",x"13",x"20",x"1A",x"F7",x"18",x"A5",x"12", -- 0x36A0
		x"69",x"28",x"85",x"12",x"90",x"02",x"E6",x"13", -- 0x36A8
		x"CA",x"D0",x"EF",x"20",x"0D",x"F7",x"A9",x"01", -- 0x36B0
		x"8D",x"68",x"02",x"AD",x"7A",x"02",x"85",x"12", -- 0x36B8
		x"AD",x"7B",x"02",x"85",x"13",x"4C",x"FE",x"F6", -- 0x36C0
		x"20",x"0D",x"F7",x"8E",x"53",x"02",x"4C",x"FE", -- 0x36C8
		x"F6",x"2A",x"2A",x"2A",x"2A",x"2A",x"2A",x"2A", -- 0x36D0
		x"2A",x"4D",x"6A",x"02",x"8D",x"6A",x"02",x"4C", -- 0x36D8
		x"FE",x"F6",x"AD",x"51",x"02",x"49",x"01",x"8D", -- 0x36E0
		x"51",x"02",x"4C",x"FE",x"F6",x"AD",x"0C",x"02", -- 0x36E8
		x"49",x"80",x"8D",x"0C",x"02",x"20",x"5A",x"F7", -- 0x36F0
		x"4C",x"FE",x"F6",x"20",x"9F",x"FA",x"AD",x"6A", -- 0x36F8
		x"02",x"0D",x"51",x"02",x"8D",x"6A",x"02",x"A9", -- 0x3700
		x"01",x"20",x"01",x"F8",x"60",x"A2",x"00",x"20", -- 0x3708
		x"DE",x"F7",x"D0",x"02",x"E8",x"E8",x"8E",x"69", -- 0x3710
		x"02",x"60",x"A0",x"27",x"A9",x"20",x"91",x"12", -- 0x3718
		x"88",x"10",x"FB",x"A0",x"00",x"AD",x"6B",x"02", -- 0x3720
		x"91",x"12",x"AD",x"6C",x"02",x"C8",x"91",x"12", -- 0x3728
		x"60",x"A0",x"00",x"8C",x"63",x"02",x"8D",x"64", -- 0x3730
		x"02",x"0A",x"2E",x"63",x"02",x"0A",x"2E",x"63", -- 0x3738
		x"02",x"18",x"6D",x"64",x"02",x"90",x"03",x"EE", -- 0x3740
		x"63",x"02",x"0A",x"2E",x"63",x"02",x"0A",x"2E", -- 0x3748
		x"63",x"02",x"0A",x"2E",x"63",x"02",x"AC",x"63", -- 0x3750
		x"02",x"60",x"AD",x"0C",x"02",x"10",x"07",x"A9", -- 0x3758
		x"70",x"A0",x"F7",x"4C",x"6A",x"F7",x"A9",x"76", -- 0x3760
		x"A0",x"F7",x"A2",x"23",x"20",x"65",x"F8",x"60", -- 0x3768
		x"07",x"43",x"41",x"50",x"53",x"00",x"07",x"20", -- 0x3770
		x"20",x"20",x"20",x"00",x"48",x"08",x"98",x"48", -- 0x3778
		x"8A",x"48",x"D8",x"E0",x"13",x"F0",x"46",x"E0", -- 0x3780
		x"14",x"F0",x"42",x"E0",x"06",x"F0",x"3E",x"AD", -- 0x3788
		x"6A",x"02",x"29",x"02",x"F0",x"3A",x"8A",x"C9", -- 0x3790
		x"20",x"90",x"32",x"AD",x"6A",x"02",x"29",x"10", -- 0x3798
		x"F0",x"13",x"8A",x"38",x"E9",x"40",x"30",x"09", -- 0x37A0
		x"29",x"1F",x"20",x"E4",x"F7",x"A9",x"1B",x"D0", -- 0x37A8
		x"1C",x"A9",x"20",x"10",x"F5",x"E0",x"7F",x"F0", -- 0x37B0
		x"08",x"68",x"48",x"20",x"E4",x"F7",x"4C",x"D0", -- 0x37B8
		x"F7",x"A9",x"08",x"20",x"02",x"F6",x"A9",x"20", -- 0x37C0
		x"20",x"E4",x"F7",x"A9",x"08",x"20",x"02",x"F6", -- 0x37C8
		x"68",x"AA",x"68",x"A8",x"28",x"68",x"60",x"AD", -- 0x37D0
		x"69",x"02",x"29",x"FE",x"D0",x"05",x"AD",x"6A", -- 0x37D8
		x"02",x"29",x"20",x"60",x"48",x"AC",x"69",x"02", -- 0x37E0
		x"91",x"12",x"2C",x"6A",x"02",x"50",x"0B",x"AD", -- 0x37E8
		x"69",x"02",x"18",x"69",x"28",x"A8",x"68",x"48", -- 0x37F0
		x"91",x"12",x"A9",x"09",x"20",x"02",x"F6",x"68", -- 0x37F8
		x"60",x"2D",x"6A",x"02",x"4A",x"6A",x"8D",x"65", -- 0x3800
		x"02",x"AC",x"69",x"02",x"B1",x"12",x"29",x"7F", -- 0x3808
		x"0D",x"65",x"02",x"91",x"12",x"60",x"A9",x"00", -- 0x3810
		x"85",x"0C",x"A9",x"B9",x"85",x"0D",x"A9",x"00", -- 0x3818
		x"20",x"2D",x"F8",x"A0",x"BA",x"84",x"0D",x"A9", -- 0x3820
		x"20",x"20",x"2D",x"F8",x"60",x"A0",x"00",x"48", -- 0x3828
		x"20",x"54",x"F8",x"91",x"0C",x"C8",x"68",x"48", -- 0x3830
		x"20",x"52",x"F8",x"68",x"48",x"20",x"50",x"F8", -- 0x3838
		x"91",x"0C",x"C8",x"C0",x"00",x"F0",x"07",x"68", -- 0x3840
		x"18",x"69",x"01",x"4C",x"2F",x"F8",x"68",x"60", -- 0x3848
		x"4A",x"4A",x"4A",x"4A",x"29",x"03",x"AA",x"BD", -- 0x3850
		x"61",x"F8",x"91",x"0C",x"C8",x"91",x"0C",x"C8", -- 0x3858
		x"60",x"00",x"38",x"07",x"3F",x"85",x"0C",x"84", -- 0x3860
		x"0D",x"AD",x"1F",x"02",x"D0",x"0D",x"A0",x"00", -- 0x3868
		x"B1",x"0C",x"F0",x"07",x"9D",x"80",x"BB",x"E8", -- 0x3870
		x"C8",x"D0",x"F5",x"60",x"4C",x"7C",x"F7",x"4C", -- 0x3878
		x"78",x"EB",x"4C",x"C1",x"F5",x"4C",x"65",x"F8", -- 0x3880
		x"4C",x"22",x"EE",x"4C",x"B2",x"F8",x"40",x"A2", -- 0x3888
		x"FF",x"9A",x"58",x"D8",x"A2",x"12",x"BD",x"7C", -- 0x3890
		x"F8",x"9D",x"38",x"02",x"CA",x"10",x"F7",x"A9", -- 0x3898
		x"20",x"8D",x"4E",x"02",x"A9",x"04",x"8D",x"4F", -- 0x38A0
		x"02",x"20",x"14",x"FA",x"20",x"B8",x"F8",x"4C", -- 0x38A8
		x"CC",x"EC",x"20",x"B8",x"F8",x"4C",x"71",x"C4", -- 0x38B0
		x"20",x"AA",x"F9",x"A9",x"07",x"A2",x"40",x"20", -- 0x38B8
		x"90",x"F5",x"20",x"E0",x"ED",x"20",x"0E",x"F9", -- 0x38C0
		x"A9",x"FF",x"8D",x"0C",x"02",x"20",x"C9",x"F9", -- 0x38C8
		x"A2",x"05",x"20",x"82",x"F9",x"20",x"16",x"F8", -- 0x38D0
		x"20",x"5A",x"F7",x"60",x"48",x"8A",x"48",x"A9", -- 0x38D8
		x"01",x"8D",x"1F",x"02",x"A9",x"BF",x"8D",x"7B", -- 0x38E0
		x"02",x"8D",x"79",x"02",x"A9",x"68",x"8D",x"7A", -- 0x38E8
		x"02",x"A9",x"90",x"8D",x"78",x"02",x"A9",x"03", -- 0x38F0
		x"8D",x"7E",x"02",x"A9",x"00",x"8D",x"7D",x"02", -- 0x38F8
		x"A9",x"50",x"8D",x"7C",x"02",x"A2",x"0C",x"20", -- 0x3900
		x"38",x"02",x"68",x"AA",x"68",x"60",x"48",x"A9", -- 0x3908
		x"03",x"8D",x"6A",x"02",x"A9",x"00",x"8D",x"6C", -- 0x3910
		x"02",x"A9",x"17",x"8D",x"6B",x"02",x"68",x"60", -- 0x3918
		x"48",x"AD",x"1F",x"02",x"D0",x"05",x"A2",x"0B", -- 0x3920
		x"20",x"82",x"F9",x"A9",x"FE",x"2D",x"6A",x"02", -- 0x3928
		x"8D",x"6A",x"02",x"A9",x"1E",x"8D",x"DF",x"BF", -- 0x3930
		x"A9",x"40",x"8D",x"00",x"A0",x"A2",x"17",x"20", -- 0x3938
		x"82",x"F9",x"A9",x"00",x"8D",x"19",x"02",x"8D", -- 0x3940
		x"1A",x"02",x"85",x"10",x"A9",x"A0",x"85",x"11", -- 0x3948
		x"A9",x"20",x"8D",x"15",x"02",x"A9",x"FF",x"8D", -- 0x3950
		x"13",x"02",x"20",x"DC",x"F8",x"A9",x"01",x"0D", -- 0x3958
		x"6A",x"02",x"8D",x"6A",x"02",x"68",x"60",x"48", -- 0x3960
		x"A9",x"FE",x"2D",x"6A",x"02",x"8D",x"6A",x"02", -- 0x3968
		x"A2",x"11",x"20",x"82",x"F9",x"20",x"C9",x"F9", -- 0x3970
		x"A9",x"01",x"0D",x"6A",x"02",x"8D",x"6A",x"02", -- 0x3978
		x"68",x"60",x"A0",x"06",x"BD",x"92",x"F9",x"99", -- 0x3980
		x"0B",x"00",x"CA",x"88",x"D0",x"F6",x"20",x"C4", -- 0x3988
		x"ED",x"60",x"78",x"FC",x"00",x"B5",x"00",x"03", -- 0x3990
		x"00",x"B4",x"00",x"98",x"80",x"07",x"00",x"98", -- 0x3998
		x"00",x"B4",x"80",x"07",x"00",x"A0",x"01",x"A0", -- 0x39A0
		x"3F",x"1F",x"A9",x"FF",x"8D",x"03",x"03",x"A9", -- 0x39A8
		x"F7",x"8D",x"02",x"03",x"A9",x"B7",x"8D",x"00", -- 0x39B0
		x"03",x"A9",x"DD",x"8D",x"0C",x"03",x"A9",x"7F", -- 0x39B8
		x"8D",x"0E",x"03",x"A9",x"00",x"8D",x"0B",x"03", -- 0x39C0
		x"60",x"A9",x"1A",x"20",x"07",x"FA",x"A9",x"20", -- 0x39C8
		x"A0",x"28",x"99",x"7F",x"BB",x"88",x"D0",x"FA", -- 0x39D0
		x"A9",x"00",x"8D",x"1F",x"02",x"A9",x"BB",x"8D", -- 0x39D8
		x"7B",x"02",x"8D",x"79",x"02",x"A9",x"A8",x"8D", -- 0x39E0
		x"7A",x"02",x"A9",x"D0",x"8D",x"78",x"02",x"A9", -- 0x39E8
		x"1B",x"8D",x"7E",x"02",x"A9",x"04",x"8D",x"7D", -- 0x39F0
		x"02",x"A9",x"10",x"8D",x"7C",x"02",x"A2",x"0C", -- 0x39F8
		x"20",x"38",x"02",x"20",x"5A",x"F7",x"60",x"8D", -- 0x3A00
		x"DF",x"BF",x"A9",x"02",x"A2",x"00",x"A0",x"03", -- 0x3A08
		x"20",x"C9",x"EE",x"60",x"A0",x"00",x"8C",x"60", -- 0x3A10
		x"02",x"8C",x"20",x"02",x"8C",x"00",x"05",x"84", -- 0x3A18
		x"0E",x"88",x"84",x"0C",x"8C",x"00",x"45",x"AD", -- 0x3A20
		x"00",x"05",x"D0",x"04",x"A9",x"C0",x"D0",x"05", -- 0x3A28
		x"EE",x"20",x"02",x"A9",x"40",x"85",x"0F",x"C8", -- 0x3A30
		x"A9",x"03",x"85",x"0D",x"E6",x"0C",x"D0",x"02", -- 0x3A38
--		x"A9",x"BF",x"85",x"0D",x"E6",x"0C",x"D0",x"02", -- 0x3A38 -- To speed up simulation
		x"E6",x"0D",x"A5",x"0C",x"C5",x"0E",x"D0",x"06", -- 0x3A40
		x"A5",x"0D",x"C5",x"0F",x"F0",x"0F",x"A9",x"AA", -- 0x3A48
		x"91",x"0C",x"D1",x"0C",x"D0",x"07",x"4A",x"91", -- 0x3A50
		x"0C",x"D1",x"0C",x"F0",x"DF",x"38",x"A5",x"0F", -- 0x3A58
		x"E9",x"28",x"85",x"0F",x"A5",x"0E",x"C5",x"0C", -- 0x3A60
		x"A5",x"0F",x"E5",x"0D",x"90",x"09",x"A5",x"0C", -- 0x3A68
		x"A4",x"0D",x"EE",x"60",x"02",x"D0",x"04",x"A5", -- 0x3A70
		x"0E",x"A4",x"0F",x"85",x"A6",x"84",x"A7",x"8D", -- 0x3A78
		x"C1",x"02",x"8C",x"C2",x"02",x"60",x"08",x"78", -- 0x3A80
		x"86",x"14",x"84",x"15",x"A0",x"00",x"B1",x"14", -- 0x3A88
		x"AA",x"98",x"48",x"20",x"90",x"F5",x"68",x"A8", -- 0x3A90
		x"C8",x"C0",x"0E",x"D0",x"F1",x"28",x"60",x"A2", -- 0x3A98
		x"A7",x"A0",x"FA",x"20",x"86",x"FA",x"60",x"18", -- 0x3AA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"10", -- 0x3AA8
		x"00",x"00",x"00",x"0F",x"00",x"A2",x"BD",x"A0", -- 0x3AB0
		x"FA",x"20",x"86",x"FA",x"60",x"00",x"00",x"00", -- 0x3AB8
		x"00",x"00",x"00",x"0F",x"07",x"10",x"10",x"10", -- 0x3AC0
		x"00",x"08",x"00",x"A2",x"D3",x"A0",x"FA",x"20", -- 0x3AC8
		x"86",x"FA",x"60",x"00",x"00",x"00",x"00",x"00", -- 0x3AD0
		x"00",x"1F",x"07",x"10",x"10",x"10",x"00",x"18", -- 0x3AD8
		x"00",x"A2",x"06",x"A0",x"FB",x"20",x"86",x"FA", -- 0x3AE0
		x"A9",x"00",x"AA",x"8A",x"48",x"A9",x"00",x"20", -- 0x3AE8
		x"90",x"F5",x"A2",x"00",x"CA",x"D0",x"FD",x"68", -- 0x3AF0
		x"AA",x"E8",x"E0",x"70",x"D0",x"ED",x"A9",x"08", -- 0x3AF8
		x"A2",x"00",x"20",x"90",x"F5",x"60",x"00",x"00", -- 0x3B00
		x"00",x"00",x"00",x"00",x"00",x"3E",x"0F",x"00", -- 0x3B08
		x"00",x"00",x"00",x"00",x"A2",x"1C",x"A0",x"FB", -- 0x3B10
		x"20",x"86",x"FA",x"60",x"1F",x"00",x"00",x"00", -- 0x3B18
		x"00",x"00",x"00",x"3E",x"10",x"00",x"00",x"1F", -- 0x3B20
		x"00",x"00",x"A2",x"32",x"A0",x"FB",x"20",x"86", -- 0x3B28
		x"FA",x"60",x"2F",x"00",x"00",x"00",x"00",x"00", -- 0x3B30
		x"00",x"3E",x"10",x"00",x"00",x"1F",x"00",x"00", -- 0x3B38
		x"AD",x"E1",x"02",x"C9",x"01",x"D0",x"22",x"A9", -- 0x3B40
		x"00",x"AE",x"E3",x"02",x"20",x"90",x"F5",x"A9", -- 0x3B48
		x"01",x"AE",x"E4",x"02",x"20",x"90",x"F5",x"AD", -- 0x3B50
		x"E5",x"02",x"29",x"0F",x"D0",x"04",x"A2",x"10", -- 0x3B58
		x"D0",x"01",x"AA",x"A9",x"08",x"20",x"90",x"F5", -- 0x3B60
		x"60",x"C9",x"02",x"D0",x"22",x"A9",x"02",x"AE", -- 0x3B68
		x"E3",x"02",x"20",x"90",x"F5",x"A9",x"03",x"AE", -- 0x3B70
		x"E4",x"02",x"20",x"90",x"F5",x"AD",x"E5",x"02", -- 0x3B78
		x"29",x"0F",x"D0",x"04",x"A2",x"10",x"D0",x"01", -- 0x3B80
		x"AA",x"A9",x"09",x"20",x"90",x"F5",x"60",x"C9", -- 0x3B88
		x"03",x"D0",x"22",x"A9",x"04",x"AE",x"E3",x"02", -- 0x3B90
		x"20",x"90",x"F5",x"A9",x"05",x"AE",x"E4",x"02", -- 0x3B98
		x"20",x"90",x"F5",x"AD",x"E5",x"02",x"29",x"0F", -- 0x3BA0
		x"D0",x"04",x"A2",x"10",x"D0",x"01",x"AA",x"A9", -- 0x3BA8
		x"0A",x"20",x"90",x"F5",x"60",x"A9",x"06",x"AE", -- 0x3BB0
		x"E3",x"02",x"20",x"90",x"F5",x"AD",x"E1",x"02", -- 0x3BB8
		x"C9",x"04",x"F0",x"93",x"C9",x"05",x"F0",x"B5", -- 0x3BC0
		x"C9",x"06",x"F0",x"D7",x"EE",x"E0",x"02",x"60", -- 0x3BC8
		x"AD",x"E3",x"02",x"0A",x"0A",x"0A",x"0D",x"E1", -- 0x3BD0
		x"02",x"49",x"3F",x"AA",x"A9",x"07",x"20",x"90", -- 0x3BD8
		x"F5",x"18",x"AD",x"E7",x"02",x"0A",x"8D",x"E7", -- 0x3BE0
		x"02",x"AD",x"E8",x"02",x"2A",x"8D",x"E8",x"02", -- 0x3BE8
		x"A9",x"0B",x"AE",x"E7",x"02",x"20",x"90",x"F5", -- 0x3BF0
		x"A9",x"0C",x"AE",x"E8",x"02",x"20",x"90",x"F5", -- 0x3BF8
		x"AD",x"E5",x"02",x"29",x"07",x"A8",x"B9",x"10", -- 0x3C00
		x"FC",x"AA",x"A9",x"0D",x"20",x"90",x"F5",x"60", -- 0x3C08
		x"00",x"00",x"04",x"08",x"0A",x"0B",x"0C",x"0D", -- 0x3C10
		x"A2",x"E1",x"A9",x"04",x"20",x"E4",x"F2",x"B0", -- 0x3C18
		x"39",x"A2",x"E3",x"A9",x"08",x"20",x"F8",x"F2", -- 0x3C20
		x"B0",x"30",x"A2",x"E5",x"A9",x"0D",x"20",x"E4", -- 0x3C28
		x"F2",x"B0",x"27",x"AC",x"E3",x"02",x"AE",x"E5", -- 0x3C30
		x"02",x"BD",x"5E",x"FC",x"8D",x"E4",x"02",x"BD", -- 0x3C38
		x"6B",x"FC",x"8D",x"E3",x"02",x"AD",x"E7",x"02", -- 0x3C40
		x"8D",x"E5",x"02",x"88",x"30",x"09",x"4E",x"E4", -- 0x3C48
		x"02",x"6E",x"E3",x"02",x"4C",x"4B",x"FC",x"4C", -- 0x3C50
		x"40",x"FB",x"EE",x"E0",x"02",x"60",x"00",x"07", -- 0x3C58
		x"07",x"06",x"06",x"05",x"05",x"05",x"04",x"04", -- 0x3C60
		x"04",x"04",x"03",x"00",x"77",x"0B",x"A6",x"47", -- 0x3C68
		x"EC",x"97",x"47",x"FB",x"B3",x"70",x"30",x"F4", -- 0x3C70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C78
		x"08",x"08",x"08",x"08",x"08",x"00",x"08",x"00", -- 0x3C80
		x"14",x"14",x"14",x"00",x"00",x"00",x"00",x"00", -- 0x3C88
		x"14",x"14",x"3E",x"14",x"3E",x"14",x"14",x"00", -- 0x3C90
		x"08",x"1E",x"28",x"1C",x"0A",x"3C",x"08",x"00", -- 0x3C98
		x"30",x"32",x"04",x"08",x"10",x"26",x"06",x"00", -- 0x3CA0
		x"10",x"28",x"28",x"10",x"2A",x"24",x"1A",x"00", -- 0x3CA8
		x"08",x"08",x"08",x"00",x"00",x"00",x"00",x"00", -- 0x3CB0
		x"08",x"10",x"20",x"20",x"20",x"10",x"08",x"00", -- 0x3CB8
		x"08",x"04",x"02",x"02",x"02",x"04",x"08",x"00", -- 0x3CC0
		x"08",x"2A",x"1C",x"08",x"1C",x"2A",x"08",x"00", -- 0x3CC8
		x"00",x"08",x"08",x"3E",x"08",x"08",x"00",x"00", -- 0x3CD0
		x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"10", -- 0x3CD8
		x"00",x"00",x"00",x"3E",x"00",x"00",x"00",x"00", -- 0x3CE0
		x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00", -- 0x3CE8
		x"00",x"02",x"04",x"08",x"10",x"20",x"00",x"00", -- 0x3CF0
		x"1C",x"22",x"26",x"2A",x"32",x"22",x"1C",x"00", -- 0x3CF8
		x"08",x"18",x"08",x"08",x"08",x"08",x"1C",x"00", -- 0x3D00
		x"1C",x"22",x"02",x"04",x"08",x"10",x"3E",x"00", -- 0x3D08
		x"3E",x"02",x"04",x"0C",x"02",x"22",x"1C",x"00", -- 0x3D10
		x"04",x"0C",x"14",x"24",x"3E",x"04",x"04",x"00", -- 0x3D18
		x"3E",x"20",x"3C",x"02",x"02",x"22",x"1C",x"00", -- 0x3D20
		x"0C",x"10",x"20",x"3C",x"22",x"22",x"1C",x"00", -- 0x3D28
		x"3E",x"02",x"04",x"08",x"10",x"10",x"10",x"00", -- 0x3D30
		x"1C",x"22",x"22",x"1C",x"22",x"22",x"1C",x"00", -- 0x3D38
		x"1C",x"22",x"22",x"1E",x"02",x"04",x"18",x"00", -- 0x3D40
		x"00",x"00",x"08",x"00",x"00",x"08",x"00",x"00", -- 0x3D48
		x"00",x"00",x"08",x"00",x"00",x"08",x"08",x"10", -- 0x3D50
		x"04",x"08",x"10",x"20",x"10",x"08",x"04",x"00", -- 0x3D58
		x"00",x"00",x"3E",x"00",x"3E",x"00",x"00",x"00", -- 0x3D60
		x"10",x"08",x"04",x"02",x"04",x"08",x"10",x"00", -- 0x3D68
		x"1C",x"22",x"04",x"08",x"08",x"00",x"08",x"00", -- 0x3D70
		x"1C",x"22",x"2A",x"2E",x"2C",x"20",x"1E",x"00", -- 0x3D78
		x"08",x"14",x"22",x"22",x"3E",x"22",x"22",x"00", -- 0x3D80
		x"3C",x"22",x"22",x"3C",x"22",x"22",x"3C",x"00", -- 0x3D88
		x"1C",x"22",x"20",x"20",x"20",x"22",x"1C",x"00", -- 0x3D90
		x"3C",x"22",x"22",x"22",x"22",x"22",x"3C",x"00", -- 0x3D98
		x"3E",x"20",x"20",x"3C",x"20",x"20",x"3E",x"00", -- 0x3DA0
		x"3E",x"20",x"20",x"3C",x"20",x"20",x"20",x"00", -- 0x3DA8
		x"1E",x"20",x"20",x"20",x"26",x"22",x"1E",x"00", -- 0x3DB0
		x"22",x"22",x"22",x"3E",x"22",x"22",x"22",x"00", -- 0x3DB8
		x"1C",x"08",x"08",x"08",x"08",x"08",x"1C",x"00", -- 0x3DC0
		x"02",x"02",x"02",x"02",x"02",x"22",x"1C",x"00", -- 0x3DC8
		x"22",x"24",x"28",x"30",x"28",x"24",x"22",x"00", -- 0x3DD0
		x"20",x"20",x"20",x"20",x"20",x"20",x"3E",x"00", -- 0x3DD8
		x"22",x"36",x"2A",x"2A",x"22",x"22",x"22",x"00", -- 0x3DE0
		x"22",x"22",x"32",x"2A",x"26",x"22",x"22",x"00", -- 0x3DE8
		x"1C",x"22",x"22",x"22",x"22",x"22",x"1C",x"00", -- 0x3DF0
		x"3C",x"22",x"22",x"3C",x"20",x"20",x"20",x"00", -- 0x3DF8
		x"1C",x"22",x"22",x"22",x"2A",x"24",x"1A",x"00", -- 0x3E00
		x"3C",x"22",x"22",x"3C",x"28",x"24",x"22",x"00", -- 0x3E08
		x"1C",x"22",x"20",x"1C",x"02",x"22",x"1C",x"00", -- 0x3E10
		x"3E",x"08",x"08",x"08",x"08",x"08",x"08",x"00", -- 0x3E18
		x"22",x"22",x"22",x"22",x"22",x"22",x"1C",x"00", -- 0x3E20
		x"22",x"22",x"22",x"22",x"22",x"14",x"08",x"00", -- 0x3E28
		x"22",x"22",x"22",x"2A",x"2A",x"36",x"22",x"00", -- 0x3E30
		x"22",x"22",x"14",x"08",x"14",x"22",x"22",x"00", -- 0x3E38
		x"22",x"22",x"14",x"08",x"08",x"08",x"08",x"00", -- 0x3E40
		x"3E",x"02",x"04",x"08",x"10",x"20",x"3E",x"00", -- 0x3E48
		x"1E",x"10",x"10",x"10",x"10",x"10",x"1E",x"00", -- 0x3E50
		x"00",x"20",x"10",x"08",x"04",x"02",x"00",x"00", -- 0x3E58
		x"3C",x"04",x"04",x"04",x"04",x"04",x"3C",x"00", -- 0x3E60
		x"08",x"14",x"2A",x"08",x"08",x"08",x"08",x"00", -- 0x3E68
		x"0E",x"10",x"10",x"10",x"3C",x"10",x"3E",x"00", -- 0x3E70
		x"0C",x"12",x"2D",x"29",x"29",x"2D",x"12",x"0C", -- 0x3E78
		x"00",x"00",x"1C",x"02",x"1E",x"22",x"1E",x"00", -- 0x3E80
		x"20",x"20",x"3C",x"22",x"22",x"22",x"3C",x"00", -- 0x3E88
		x"00",x"00",x"1E",x"20",x"20",x"20",x"1E",x"00", -- 0x3E90
		x"02",x"02",x"1E",x"22",x"22",x"22",x"1E",x"00", -- 0x3E98
		x"00",x"00",x"1C",x"22",x"3E",x"20",x"1E",x"00", -- 0x3EA0
		x"0C",x"12",x"10",x"3C",x"10",x"10",x"10",x"00", -- 0x3EA8
		x"00",x"00",x"1C",x"22",x"22",x"1E",x"02",x"1C", -- 0x3EB0
		x"20",x"20",x"3C",x"22",x"22",x"22",x"22",x"00", -- 0x3EB8
		x"08",x"00",x"18",x"08",x"08",x"08",x"1C",x"00", -- 0x3EC0
		x"04",x"00",x"0C",x"04",x"04",x"04",x"24",x"18", -- 0x3EC8
		x"20",x"20",x"22",x"24",x"38",x"24",x"22",x"00", -- 0x3ED0
		x"18",x"08",x"08",x"08",x"08",x"08",x"1C",x"00", -- 0x3ED8
		x"00",x"00",x"36",x"2A",x"2A",x"2A",x"22",x"00", -- 0x3EE0
		x"00",x"00",x"3C",x"22",x"22",x"22",x"22",x"00", -- 0x3EE8
		x"00",x"00",x"1C",x"22",x"22",x"22",x"1C",x"00", -- 0x3EF0
		x"00",x"00",x"3C",x"22",x"22",x"3C",x"20",x"20", -- 0x3EF8
		x"00",x"00",x"1E",x"22",x"22",x"1E",x"02",x"02", -- 0x3F00
		x"00",x"00",x"2E",x"30",x"20",x"20",x"20",x"00", -- 0x3F08
		x"00",x"00",x"1E",x"20",x"1C",x"02",x"3C",x"00", -- 0x3F10
		x"10",x"10",x"3C",x"10",x"10",x"12",x"0C",x"00", -- 0x3F18
		x"00",x"00",x"22",x"22",x"22",x"26",x"1A",x"00", -- 0x3F20
		x"00",x"00",x"22",x"22",x"22",x"14",x"08",x"00", -- 0x3F28
		x"00",x"00",x"22",x"22",x"2A",x"2A",x"36",x"00", -- 0x3F30
		x"00",x"00",x"22",x"14",x"08",x"14",x"22",x"00", -- 0x3F38
		x"00",x"00",x"22",x"22",x"22",x"1E",x"02",x"1C", -- 0x3F40
		x"00",x"00",x"3E",x"04",x"08",x"10",x"3E",x"00", -- 0x3F48
		x"0E",x"18",x"18",x"30",x"18",x"18",x"0E",x"00", -- 0x3F50
		x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08", -- 0x3F58
		x"38",x"0C",x"0C",x"06",x"0C",x"0C",x"38",x"00", -- 0x3F60
		x"2A",x"15",x"2A",x"15",x"2A",x"15",x"2A",x"15", -- 0x3F68
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F", -- 0x3F70
		x"37",x"EA",x"ED",x"EB",x"20",x"F5",x"F9",x"38", -- 0x3F78
		x"EE",x"F4",x"36",x"39",x"2C",x"E9",x"E8",x"EC", -- 0x3F80
		x"35",x"F2",x"E2",x"3B",x"2E",x"EF",x"E7",x"30", -- 0x3F88
		x"F6",x"E6",x"34",x"2D",x"0B",x"F0",x"E5",x"2F", -- 0x3F90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F98
		x"31",x"1B",x"FA",x"00",x"08",x"7F",x"E1",x"0D", -- 0x3FA0
		x"F8",x"F1",x"32",x"5C",x"0A",x"5D",x"F3",x"00", -- 0x3FA8
		x"33",x"E4",x"E3",x"27",x"09",x"5B",x"F7",x"3D", -- 0x3FB0
		x"26",x"4A",x"4D",x"4B",x"20",x"55",x"59",x"2A", -- 0x3FB8
		x"4E",x"54",x"5E",x"28",x"3C",x"49",x"48",x"4C", -- 0x3FC0
		x"25",x"52",x"42",x"3A",x"3E",x"4F",x"47",x"29", -- 0x3FC8
		x"56",x"46",x"24",x"5F",x"0B",x"50",x"45",x"3F", -- 0x3FD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FD8
		x"21",x"1B",x"5A",x"00",x"08",x"7F",x"41",x"0D", -- 0x3FE0
		x"58",x"51",x"40",x"7C",x"0A",x"7D",x"53",x"00", -- 0x3FE8
		x"23",x"44",x"43",x"22",x"09",x"7B",x"57",x"2B", -- 0x3FF0
		x"D0",x"01",x"47",x"02",x"8F",x"F8",x"44",x"02"  -- 0x3FF8
	);

begin

	p_rom : process(CLK)
	begin
		if (rising_edge(CLK)) then
			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
